`timescale 1 ns / 1 ps

(* CORE_GENERATION_INFO = "unikernel_unikernel,hls_ip_2022_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcu280-fsvh2892-2L-e,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2174,HLS_SYN_LUT=3944,HLS_VERSION=2022_2}" *)


module unikernel
(
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  ap_clk,
  ap_rst_n,
  interrupt,
  m_axi_in_0_ARADDR,
  m_axi_in_0_ARBURST,
  m_axi_in_0_ARCACHE,
  m_axi_in_0_ARID,
  m_axi_in_0_ARLEN,
  m_axi_in_0_ARLOCK,
  m_axi_in_0_ARPROT,
  m_axi_in_0_ARQOS,
  m_axi_in_0_ARREADY,
  m_axi_in_0_ARSIZE,
  m_axi_in_0_ARVALID,
  m_axi_in_0_AWADDR,
  m_axi_in_0_AWBURST,
  m_axi_in_0_AWCACHE,
  m_axi_in_0_AWID,
  m_axi_in_0_AWLEN,
  m_axi_in_0_AWLOCK,
  m_axi_in_0_AWPROT,
  m_axi_in_0_AWQOS,
  m_axi_in_0_AWREADY,
  m_axi_in_0_AWSIZE,
  m_axi_in_0_AWVALID,
  m_axi_in_0_BID,
  m_axi_in_0_BREADY,
  m_axi_in_0_BRESP,
  m_axi_in_0_BVALID,
  m_axi_in_0_RDATA,
  m_axi_in_0_RID,
  m_axi_in_0_RLAST,
  m_axi_in_0_RREADY,
  m_axi_in_0_RRESP,
  m_axi_in_0_RVALID,
  m_axi_in_0_WDATA,
  m_axi_in_0_WLAST,
  m_axi_in_0_WREADY,
  m_axi_in_0_WSTRB,
  m_axi_in_0_WVALID,
  m_axi_out_0_ARADDR,
  m_axi_out_0_ARBURST,
  m_axi_out_0_ARCACHE,
  m_axi_out_0_ARID,
  m_axi_out_0_ARLEN,
  m_axi_out_0_ARLOCK,
  m_axi_out_0_ARPROT,
  m_axi_out_0_ARQOS,
  m_axi_out_0_ARREADY,
  m_axi_out_0_ARSIZE,
  m_axi_out_0_ARVALID,
  m_axi_out_0_AWADDR,
  m_axi_out_0_AWBURST,
  m_axi_out_0_AWCACHE,
  m_axi_out_0_AWID,
  m_axi_out_0_AWLEN,
  m_axi_out_0_AWLOCK,
  m_axi_out_0_AWPROT,
  m_axi_out_0_AWQOS,
  m_axi_out_0_AWREADY,
  m_axi_out_0_AWSIZE,
  m_axi_out_0_AWVALID,
  m_axi_out_0_BID,
  m_axi_out_0_BREADY,
  m_axi_out_0_BRESP,
  m_axi_out_0_BVALID,
  m_axi_out_0_RDATA,
  m_axi_out_0_RID,
  m_axi_out_0_RLAST,
  m_axi_out_0_RREADY,
  m_axi_out_0_RRESP,
  m_axi_out_0_RVALID,
  m_axi_out_0_WDATA,
  m_axi_out_0_WLAST,
  m_axi_out_0_WREADY,
  m_axi_out_0_WSTRB,
  m_axi_out_0_WVALID,
  m_axi_in_1_ARADDR,
  m_axi_in_1_ARBURST,
  m_axi_in_1_ARCACHE,
  m_axi_in_1_ARID,
  m_axi_in_1_ARLEN,
  m_axi_in_1_ARLOCK,
  m_axi_in_1_ARPROT,
  m_axi_in_1_ARQOS,
  m_axi_in_1_ARREADY,
  m_axi_in_1_ARSIZE,
  m_axi_in_1_ARVALID,
  m_axi_in_1_AWADDR,
  m_axi_in_1_AWBURST,
  m_axi_in_1_AWCACHE,
  m_axi_in_1_AWID,
  m_axi_in_1_AWLEN,
  m_axi_in_1_AWLOCK,
  m_axi_in_1_AWPROT,
  m_axi_in_1_AWQOS,
  m_axi_in_1_AWREADY,
  m_axi_in_1_AWSIZE,
  m_axi_in_1_AWVALID,
  m_axi_in_1_BID,
  m_axi_in_1_BREADY,
  m_axi_in_1_BRESP,
  m_axi_in_1_BVALID,
  m_axi_in_1_RDATA,
  m_axi_in_1_RID,
  m_axi_in_1_RLAST,
  m_axi_in_1_RREADY,
  m_axi_in_1_RRESP,
  m_axi_in_1_RVALID,
  m_axi_in_1_WDATA,
  m_axi_in_1_WLAST,
  m_axi_in_1_WREADY,
  m_axi_in_1_WSTRB,
  m_axi_in_1_WVALID,
  m_axi_out_1_ARADDR,
  m_axi_out_1_ARBURST,
  m_axi_out_1_ARCACHE,
  m_axi_out_1_ARID,
  m_axi_out_1_ARLEN,
  m_axi_out_1_ARLOCK,
  m_axi_out_1_ARPROT,
  m_axi_out_1_ARQOS,
  m_axi_out_1_ARREADY,
  m_axi_out_1_ARSIZE,
  m_axi_out_1_ARVALID,
  m_axi_out_1_AWADDR,
  m_axi_out_1_AWBURST,
  m_axi_out_1_AWCACHE,
  m_axi_out_1_AWID,
  m_axi_out_1_AWLEN,
  m_axi_out_1_AWLOCK,
  m_axi_out_1_AWPROT,
  m_axi_out_1_AWQOS,
  m_axi_out_1_AWREADY,
  m_axi_out_1_AWSIZE,
  m_axi_out_1_AWVALID,
  m_axi_out_1_BID,
  m_axi_out_1_BREADY,
  m_axi_out_1_BRESP,
  m_axi_out_1_BVALID,
  m_axi_out_1_RDATA,
  m_axi_out_1_RID,
  m_axi_out_1_RLAST,
  m_axi_out_1_RREADY,
  m_axi_out_1_RRESP,
  m_axi_out_1_RVALID,
  m_axi_out_1_WDATA,
  m_axi_out_1_WLAST,
  m_axi_out_1_WREADY,
  m_axi_out_1_WSTRB,
  m_axi_out_1_WVALID,
  m_axi_in_2_ARADDR,
  m_axi_in_2_ARBURST,
  m_axi_in_2_ARCACHE,
  m_axi_in_2_ARID,
  m_axi_in_2_ARLEN,
  m_axi_in_2_ARLOCK,
  m_axi_in_2_ARPROT,
  m_axi_in_2_ARQOS,
  m_axi_in_2_ARREADY,
  m_axi_in_2_ARSIZE,
  m_axi_in_2_ARVALID,
  m_axi_in_2_AWADDR,
  m_axi_in_2_AWBURST,
  m_axi_in_2_AWCACHE,
  m_axi_in_2_AWID,
  m_axi_in_2_AWLEN,
  m_axi_in_2_AWLOCK,
  m_axi_in_2_AWPROT,
  m_axi_in_2_AWQOS,
  m_axi_in_2_AWREADY,
  m_axi_in_2_AWSIZE,
  m_axi_in_2_AWVALID,
  m_axi_in_2_BID,
  m_axi_in_2_BREADY,
  m_axi_in_2_BRESP,
  m_axi_in_2_BVALID,
  m_axi_in_2_RDATA,
  m_axi_in_2_RID,
  m_axi_in_2_RLAST,
  m_axi_in_2_RREADY,
  m_axi_in_2_RRESP,
  m_axi_in_2_RVALID,
  m_axi_in_2_WDATA,
  m_axi_in_2_WLAST,
  m_axi_in_2_WREADY,
  m_axi_in_2_WSTRB,
  m_axi_in_2_WVALID,
  m_axi_out_2_ARADDR,
  m_axi_out_2_ARBURST,
  m_axi_out_2_ARCACHE,
  m_axi_out_2_ARID,
  m_axi_out_2_ARLEN,
  m_axi_out_2_ARLOCK,
  m_axi_out_2_ARPROT,
  m_axi_out_2_ARQOS,
  m_axi_out_2_ARREADY,
  m_axi_out_2_ARSIZE,
  m_axi_out_2_ARVALID,
  m_axi_out_2_AWADDR,
  m_axi_out_2_AWBURST,
  m_axi_out_2_AWCACHE,
  m_axi_out_2_AWID,
  m_axi_out_2_AWLEN,
  m_axi_out_2_AWLOCK,
  m_axi_out_2_AWPROT,
  m_axi_out_2_AWQOS,
  m_axi_out_2_AWREADY,
  m_axi_out_2_AWSIZE,
  m_axi_out_2_AWVALID,
  m_axi_out_2_BID,
  m_axi_out_2_BREADY,
  m_axi_out_2_BRESP,
  m_axi_out_2_BVALID,
  m_axi_out_2_RDATA,
  m_axi_out_2_RID,
  m_axi_out_2_RLAST,
  m_axi_out_2_RREADY,
  m_axi_out_2_RRESP,
  m_axi_out_2_RVALID,
  m_axi_out_2_WDATA,
  m_axi_out_2_WLAST,
  m_axi_out_2_WREADY,
  m_axi_out_2_WSTRB,
  m_axi_out_2_WVALID,
  m_axi_in_3_ARADDR,
  m_axi_in_3_ARBURST,
  m_axi_in_3_ARCACHE,
  m_axi_in_3_ARID,
  m_axi_in_3_ARLEN,
  m_axi_in_3_ARLOCK,
  m_axi_in_3_ARPROT,
  m_axi_in_3_ARQOS,
  m_axi_in_3_ARREADY,
  m_axi_in_3_ARSIZE,
  m_axi_in_3_ARVALID,
  m_axi_in_3_AWADDR,
  m_axi_in_3_AWBURST,
  m_axi_in_3_AWCACHE,
  m_axi_in_3_AWID,
  m_axi_in_3_AWLEN,
  m_axi_in_3_AWLOCK,
  m_axi_in_3_AWPROT,
  m_axi_in_3_AWQOS,
  m_axi_in_3_AWREADY,
  m_axi_in_3_AWSIZE,
  m_axi_in_3_AWVALID,
  m_axi_in_3_BID,
  m_axi_in_3_BREADY,
  m_axi_in_3_BRESP,
  m_axi_in_3_BVALID,
  m_axi_in_3_RDATA,
  m_axi_in_3_RID,
  m_axi_in_3_RLAST,
  m_axi_in_3_RREADY,
  m_axi_in_3_RRESP,
  m_axi_in_3_RVALID,
  m_axi_in_3_WDATA,
  m_axi_in_3_WLAST,
  m_axi_in_3_WREADY,
  m_axi_in_3_WSTRB,
  m_axi_in_3_WVALID,
  m_axi_out_3_ARADDR,
  m_axi_out_3_ARBURST,
  m_axi_out_3_ARCACHE,
  m_axi_out_3_ARID,
  m_axi_out_3_ARLEN,
  m_axi_out_3_ARLOCK,
  m_axi_out_3_ARPROT,
  m_axi_out_3_ARQOS,
  m_axi_out_3_ARREADY,
  m_axi_out_3_ARSIZE,
  m_axi_out_3_ARVALID,
  m_axi_out_3_AWADDR,
  m_axi_out_3_AWBURST,
  m_axi_out_3_AWCACHE,
  m_axi_out_3_AWID,
  m_axi_out_3_AWLEN,
  m_axi_out_3_AWLOCK,
  m_axi_out_3_AWPROT,
  m_axi_out_3_AWQOS,
  m_axi_out_3_AWREADY,
  m_axi_out_3_AWSIZE,
  m_axi_out_3_AWVALID,
  m_axi_out_3_BID,
  m_axi_out_3_BREADY,
  m_axi_out_3_BRESP,
  m_axi_out_3_BVALID,
  m_axi_out_3_RDATA,
  m_axi_out_3_RID,
  m_axi_out_3_RLAST,
  m_axi_out_3_RREADY,
  m_axi_out_3_RRESP,
  m_axi_out_3_RVALID,
  m_axi_out_3_WDATA,
  m_axi_out_3_WLAST,
  m_axi_out_3_WREADY,
  m_axi_out_3_WSTRB,
  m_axi_out_3_WVALID,
  m_axi_in_4_ARADDR,
  m_axi_in_4_ARBURST,
  m_axi_in_4_ARCACHE,
  m_axi_in_4_ARID,
  m_axi_in_4_ARLEN,
  m_axi_in_4_ARLOCK,
  m_axi_in_4_ARPROT,
  m_axi_in_4_ARQOS,
  m_axi_in_4_ARREADY,
  m_axi_in_4_ARSIZE,
  m_axi_in_4_ARVALID,
  m_axi_in_4_AWADDR,
  m_axi_in_4_AWBURST,
  m_axi_in_4_AWCACHE,
  m_axi_in_4_AWID,
  m_axi_in_4_AWLEN,
  m_axi_in_4_AWLOCK,
  m_axi_in_4_AWPROT,
  m_axi_in_4_AWQOS,
  m_axi_in_4_AWREADY,
  m_axi_in_4_AWSIZE,
  m_axi_in_4_AWVALID,
  m_axi_in_4_BID,
  m_axi_in_4_BREADY,
  m_axi_in_4_BRESP,
  m_axi_in_4_BVALID,
  m_axi_in_4_RDATA,
  m_axi_in_4_RID,
  m_axi_in_4_RLAST,
  m_axi_in_4_RREADY,
  m_axi_in_4_RRESP,
  m_axi_in_4_RVALID,
  m_axi_in_4_WDATA,
  m_axi_in_4_WLAST,
  m_axi_in_4_WREADY,
  m_axi_in_4_WSTRB,
  m_axi_in_4_WVALID,
  m_axi_out_4_ARADDR,
  m_axi_out_4_ARBURST,
  m_axi_out_4_ARCACHE,
  m_axi_out_4_ARID,
  m_axi_out_4_ARLEN,
  m_axi_out_4_ARLOCK,
  m_axi_out_4_ARPROT,
  m_axi_out_4_ARQOS,
  m_axi_out_4_ARREADY,
  m_axi_out_4_ARSIZE,
  m_axi_out_4_ARVALID,
  m_axi_out_4_AWADDR,
  m_axi_out_4_AWBURST,
  m_axi_out_4_AWCACHE,
  m_axi_out_4_AWID,
  m_axi_out_4_AWLEN,
  m_axi_out_4_AWLOCK,
  m_axi_out_4_AWPROT,
  m_axi_out_4_AWQOS,
  m_axi_out_4_AWREADY,
  m_axi_out_4_AWSIZE,
  m_axi_out_4_AWVALID,
  m_axi_out_4_BID,
  m_axi_out_4_BREADY,
  m_axi_out_4_BRESP,
  m_axi_out_4_BVALID,
  m_axi_out_4_RDATA,
  m_axi_out_4_RID,
  m_axi_out_4_RLAST,
  m_axi_out_4_RREADY,
  m_axi_out_4_RRESP,
  m_axi_out_4_RVALID,
  m_axi_out_4_WDATA,
  m_axi_out_4_WLAST,
  m_axi_out_4_WREADY,
  m_axi_out_4_WSTRB,
  m_axi_out_4_WVALID,
  m_axi_in_5_ARADDR,
  m_axi_in_5_ARBURST,
  m_axi_in_5_ARCACHE,
  m_axi_in_5_ARID,
  m_axi_in_5_ARLEN,
  m_axi_in_5_ARLOCK,
  m_axi_in_5_ARPROT,
  m_axi_in_5_ARQOS,
  m_axi_in_5_ARREADY,
  m_axi_in_5_ARSIZE,
  m_axi_in_5_ARVALID,
  m_axi_in_5_AWADDR,
  m_axi_in_5_AWBURST,
  m_axi_in_5_AWCACHE,
  m_axi_in_5_AWID,
  m_axi_in_5_AWLEN,
  m_axi_in_5_AWLOCK,
  m_axi_in_5_AWPROT,
  m_axi_in_5_AWQOS,
  m_axi_in_5_AWREADY,
  m_axi_in_5_AWSIZE,
  m_axi_in_5_AWVALID,
  m_axi_in_5_BID,
  m_axi_in_5_BREADY,
  m_axi_in_5_BRESP,
  m_axi_in_5_BVALID,
  m_axi_in_5_RDATA,
  m_axi_in_5_RID,
  m_axi_in_5_RLAST,
  m_axi_in_5_RREADY,
  m_axi_in_5_RRESP,
  m_axi_in_5_RVALID,
  m_axi_in_5_WDATA,
  m_axi_in_5_WLAST,
  m_axi_in_5_WREADY,
  m_axi_in_5_WSTRB,
  m_axi_in_5_WVALID,
  m_axi_out_5_ARADDR,
  m_axi_out_5_ARBURST,
  m_axi_out_5_ARCACHE,
  m_axi_out_5_ARID,
  m_axi_out_5_ARLEN,
  m_axi_out_5_ARLOCK,
  m_axi_out_5_ARPROT,
  m_axi_out_5_ARQOS,
  m_axi_out_5_ARREADY,
  m_axi_out_5_ARSIZE,
  m_axi_out_5_ARVALID,
  m_axi_out_5_AWADDR,
  m_axi_out_5_AWBURST,
  m_axi_out_5_AWCACHE,
  m_axi_out_5_AWID,
  m_axi_out_5_AWLEN,
  m_axi_out_5_AWLOCK,
  m_axi_out_5_AWPROT,
  m_axi_out_5_AWQOS,
  m_axi_out_5_AWREADY,
  m_axi_out_5_AWSIZE,
  m_axi_out_5_AWVALID,
  m_axi_out_5_BID,
  m_axi_out_5_BREADY,
  m_axi_out_5_BRESP,
  m_axi_out_5_BVALID,
  m_axi_out_5_RDATA,
  m_axi_out_5_RID,
  m_axi_out_5_RLAST,
  m_axi_out_5_RREADY,
  m_axi_out_5_RRESP,
  m_axi_out_5_RVALID,
  m_axi_out_5_WDATA,
  m_axi_out_5_WLAST,
  m_axi_out_5_WREADY,
  m_axi_out_5_WSTRB,
  m_axi_out_5_WVALID,
  m_axi_in_6_ARADDR,
  m_axi_in_6_ARBURST,
  m_axi_in_6_ARCACHE,
  m_axi_in_6_ARID,
  m_axi_in_6_ARLEN,
  m_axi_in_6_ARLOCK,
  m_axi_in_6_ARPROT,
  m_axi_in_6_ARQOS,
  m_axi_in_6_ARREADY,
  m_axi_in_6_ARSIZE,
  m_axi_in_6_ARVALID,
  m_axi_in_6_AWADDR,
  m_axi_in_6_AWBURST,
  m_axi_in_6_AWCACHE,
  m_axi_in_6_AWID,
  m_axi_in_6_AWLEN,
  m_axi_in_6_AWLOCK,
  m_axi_in_6_AWPROT,
  m_axi_in_6_AWQOS,
  m_axi_in_6_AWREADY,
  m_axi_in_6_AWSIZE,
  m_axi_in_6_AWVALID,
  m_axi_in_6_BID,
  m_axi_in_6_BREADY,
  m_axi_in_6_BRESP,
  m_axi_in_6_BVALID,
  m_axi_in_6_RDATA,
  m_axi_in_6_RID,
  m_axi_in_6_RLAST,
  m_axi_in_6_RREADY,
  m_axi_in_6_RRESP,
  m_axi_in_6_RVALID,
  m_axi_in_6_WDATA,
  m_axi_in_6_WLAST,
  m_axi_in_6_WREADY,
  m_axi_in_6_WSTRB,
  m_axi_in_6_WVALID,
  m_axi_out_6_ARADDR,
  m_axi_out_6_ARBURST,
  m_axi_out_6_ARCACHE,
  m_axi_out_6_ARID,
  m_axi_out_6_ARLEN,
  m_axi_out_6_ARLOCK,
  m_axi_out_6_ARPROT,
  m_axi_out_6_ARQOS,
  m_axi_out_6_ARREADY,
  m_axi_out_6_ARSIZE,
  m_axi_out_6_ARVALID,
  m_axi_out_6_AWADDR,
  m_axi_out_6_AWBURST,
  m_axi_out_6_AWCACHE,
  m_axi_out_6_AWID,
  m_axi_out_6_AWLEN,
  m_axi_out_6_AWLOCK,
  m_axi_out_6_AWPROT,
  m_axi_out_6_AWQOS,
  m_axi_out_6_AWREADY,
  m_axi_out_6_AWSIZE,
  m_axi_out_6_AWVALID,
  m_axi_out_6_BID,
  m_axi_out_6_BREADY,
  m_axi_out_6_BRESP,
  m_axi_out_6_BVALID,
  m_axi_out_6_RDATA,
  m_axi_out_6_RID,
  m_axi_out_6_RLAST,
  m_axi_out_6_RREADY,
  m_axi_out_6_RRESP,
  m_axi_out_6_RVALID,
  m_axi_out_6_WDATA,
  m_axi_out_6_WLAST,
  m_axi_out_6_WREADY,
  m_axi_out_6_WSTRB,
  m_axi_out_6_WVALID,
  m_axi_in_7_ARADDR,
  m_axi_in_7_ARBURST,
  m_axi_in_7_ARCACHE,
  m_axi_in_7_ARID,
  m_axi_in_7_ARLEN,
  m_axi_in_7_ARLOCK,
  m_axi_in_7_ARPROT,
  m_axi_in_7_ARQOS,
  m_axi_in_7_ARREADY,
  m_axi_in_7_ARSIZE,
  m_axi_in_7_ARVALID,
  m_axi_in_7_AWADDR,
  m_axi_in_7_AWBURST,
  m_axi_in_7_AWCACHE,
  m_axi_in_7_AWID,
  m_axi_in_7_AWLEN,
  m_axi_in_7_AWLOCK,
  m_axi_in_7_AWPROT,
  m_axi_in_7_AWQOS,
  m_axi_in_7_AWREADY,
  m_axi_in_7_AWSIZE,
  m_axi_in_7_AWVALID,
  m_axi_in_7_BID,
  m_axi_in_7_BREADY,
  m_axi_in_7_BRESP,
  m_axi_in_7_BVALID,
  m_axi_in_7_RDATA,
  m_axi_in_7_RID,
  m_axi_in_7_RLAST,
  m_axi_in_7_RREADY,
  m_axi_in_7_RRESP,
  m_axi_in_7_RVALID,
  m_axi_in_7_WDATA,
  m_axi_in_7_WLAST,
  m_axi_in_7_WREADY,
  m_axi_in_7_WSTRB,
  m_axi_in_7_WVALID,
  m_axi_out_7_ARADDR,
  m_axi_out_7_ARBURST,
  m_axi_out_7_ARCACHE,
  m_axi_out_7_ARID,
  m_axi_out_7_ARLEN,
  m_axi_out_7_ARLOCK,
  m_axi_out_7_ARPROT,
  m_axi_out_7_ARQOS,
  m_axi_out_7_ARREADY,
  m_axi_out_7_ARSIZE,
  m_axi_out_7_ARVALID,
  m_axi_out_7_AWADDR,
  m_axi_out_7_AWBURST,
  m_axi_out_7_AWCACHE,
  m_axi_out_7_AWID,
  m_axi_out_7_AWLEN,
  m_axi_out_7_AWLOCK,
  m_axi_out_7_AWPROT,
  m_axi_out_7_AWQOS,
  m_axi_out_7_AWREADY,
  m_axi_out_7_AWSIZE,
  m_axi_out_7_AWVALID,
  m_axi_out_7_BID,
  m_axi_out_7_BREADY,
  m_axi_out_7_BRESP,
  m_axi_out_7_BVALID,
  m_axi_out_7_RDATA,
  m_axi_out_7_RID,
  m_axi_out_7_RLAST,
  m_axi_out_7_RREADY,
  m_axi_out_7_RRESP,
  m_axi_out_7_RVALID,
  m_axi_out_7_WDATA,
  m_axi_out_7_WLAST,
  m_axi_out_7_WREADY,
  m_axi_out_7_WSTRB,
  m_axi_out_7_WVALID,
  m_axi_in_8_ARADDR,
  m_axi_in_8_ARBURST,
  m_axi_in_8_ARCACHE,
  m_axi_in_8_ARID,
  m_axi_in_8_ARLEN,
  m_axi_in_8_ARLOCK,
  m_axi_in_8_ARPROT,
  m_axi_in_8_ARQOS,
  m_axi_in_8_ARREADY,
  m_axi_in_8_ARSIZE,
  m_axi_in_8_ARVALID,
  m_axi_in_8_AWADDR,
  m_axi_in_8_AWBURST,
  m_axi_in_8_AWCACHE,
  m_axi_in_8_AWID,
  m_axi_in_8_AWLEN,
  m_axi_in_8_AWLOCK,
  m_axi_in_8_AWPROT,
  m_axi_in_8_AWQOS,
  m_axi_in_8_AWREADY,
  m_axi_in_8_AWSIZE,
  m_axi_in_8_AWVALID,
  m_axi_in_8_BID,
  m_axi_in_8_BREADY,
  m_axi_in_8_BRESP,
  m_axi_in_8_BVALID,
  m_axi_in_8_RDATA,
  m_axi_in_8_RID,
  m_axi_in_8_RLAST,
  m_axi_in_8_RREADY,
  m_axi_in_8_RRESP,
  m_axi_in_8_RVALID,
  m_axi_in_8_WDATA,
  m_axi_in_8_WLAST,
  m_axi_in_8_WREADY,
  m_axi_in_8_WSTRB,
  m_axi_in_8_WVALID,
  m_axi_out_8_ARADDR,
  m_axi_out_8_ARBURST,
  m_axi_out_8_ARCACHE,
  m_axi_out_8_ARID,
  m_axi_out_8_ARLEN,
  m_axi_out_8_ARLOCK,
  m_axi_out_8_ARPROT,
  m_axi_out_8_ARQOS,
  m_axi_out_8_ARREADY,
  m_axi_out_8_ARSIZE,
  m_axi_out_8_ARVALID,
  m_axi_out_8_AWADDR,
  m_axi_out_8_AWBURST,
  m_axi_out_8_AWCACHE,
  m_axi_out_8_AWID,
  m_axi_out_8_AWLEN,
  m_axi_out_8_AWLOCK,
  m_axi_out_8_AWPROT,
  m_axi_out_8_AWQOS,
  m_axi_out_8_AWREADY,
  m_axi_out_8_AWSIZE,
  m_axi_out_8_AWVALID,
  m_axi_out_8_BID,
  m_axi_out_8_BREADY,
  m_axi_out_8_BRESP,
  m_axi_out_8_BVALID,
  m_axi_out_8_RDATA,
  m_axi_out_8_RID,
  m_axi_out_8_RLAST,
  m_axi_out_8_RREADY,
  m_axi_out_8_RRESP,
  m_axi_out_8_RVALID,
  m_axi_out_8_WDATA,
  m_axi_out_8_WLAST,
  m_axi_out_8_WREADY,
  m_axi_out_8_WSTRB,
  m_axi_out_8_WVALID,
  m_axi_in_9_ARADDR,
  m_axi_in_9_ARBURST,
  m_axi_in_9_ARCACHE,
  m_axi_in_9_ARID,
  m_axi_in_9_ARLEN,
  m_axi_in_9_ARLOCK,
  m_axi_in_9_ARPROT,
  m_axi_in_9_ARQOS,
  m_axi_in_9_ARREADY,
  m_axi_in_9_ARSIZE,
  m_axi_in_9_ARVALID,
  m_axi_in_9_AWADDR,
  m_axi_in_9_AWBURST,
  m_axi_in_9_AWCACHE,
  m_axi_in_9_AWID,
  m_axi_in_9_AWLEN,
  m_axi_in_9_AWLOCK,
  m_axi_in_9_AWPROT,
  m_axi_in_9_AWQOS,
  m_axi_in_9_AWREADY,
  m_axi_in_9_AWSIZE,
  m_axi_in_9_AWVALID,
  m_axi_in_9_BID,
  m_axi_in_9_BREADY,
  m_axi_in_9_BRESP,
  m_axi_in_9_BVALID,
  m_axi_in_9_RDATA,
  m_axi_in_9_RID,
  m_axi_in_9_RLAST,
  m_axi_in_9_RREADY,
  m_axi_in_9_RRESP,
  m_axi_in_9_RVALID,
  m_axi_in_9_WDATA,
  m_axi_in_9_WLAST,
  m_axi_in_9_WREADY,
  m_axi_in_9_WSTRB,
  m_axi_in_9_WVALID,
  m_axi_out_9_ARADDR,
  m_axi_out_9_ARBURST,
  m_axi_out_9_ARCACHE,
  m_axi_out_9_ARID,
  m_axi_out_9_ARLEN,
  m_axi_out_9_ARLOCK,
  m_axi_out_9_ARPROT,
  m_axi_out_9_ARQOS,
  m_axi_out_9_ARREADY,
  m_axi_out_9_ARSIZE,
  m_axi_out_9_ARVALID,
  m_axi_out_9_AWADDR,
  m_axi_out_9_AWBURST,
  m_axi_out_9_AWCACHE,
  m_axi_out_9_AWID,
  m_axi_out_9_AWLEN,
  m_axi_out_9_AWLOCK,
  m_axi_out_9_AWPROT,
  m_axi_out_9_AWQOS,
  m_axi_out_9_AWREADY,
  m_axi_out_9_AWSIZE,
  m_axi_out_9_AWVALID,
  m_axi_out_9_BID,
  m_axi_out_9_BREADY,
  m_axi_out_9_BRESP,
  m_axi_out_9_BVALID,
  m_axi_out_9_RDATA,
  m_axi_out_9_RID,
  m_axi_out_9_RLAST,
  m_axi_out_9_RREADY,
  m_axi_out_9_RRESP,
  m_axi_out_9_RVALID,
  m_axi_out_9_WDATA,
  m_axi_out_9_WLAST,
  m_axi_out_9_WREADY,
  m_axi_out_9_WSTRB,
  m_axi_out_9_WVALID,
  m_axi_in_10_ARADDR,
  m_axi_in_10_ARBURST,
  m_axi_in_10_ARCACHE,
  m_axi_in_10_ARID,
  m_axi_in_10_ARLEN,
  m_axi_in_10_ARLOCK,
  m_axi_in_10_ARPROT,
  m_axi_in_10_ARQOS,
  m_axi_in_10_ARREADY,
  m_axi_in_10_ARSIZE,
  m_axi_in_10_ARVALID,
  m_axi_in_10_AWADDR,
  m_axi_in_10_AWBURST,
  m_axi_in_10_AWCACHE,
  m_axi_in_10_AWID,
  m_axi_in_10_AWLEN,
  m_axi_in_10_AWLOCK,
  m_axi_in_10_AWPROT,
  m_axi_in_10_AWQOS,
  m_axi_in_10_AWREADY,
  m_axi_in_10_AWSIZE,
  m_axi_in_10_AWVALID,
  m_axi_in_10_BID,
  m_axi_in_10_BREADY,
  m_axi_in_10_BRESP,
  m_axi_in_10_BVALID,
  m_axi_in_10_RDATA,
  m_axi_in_10_RID,
  m_axi_in_10_RLAST,
  m_axi_in_10_RREADY,
  m_axi_in_10_RRESP,
  m_axi_in_10_RVALID,
  m_axi_in_10_WDATA,
  m_axi_in_10_WLAST,
  m_axi_in_10_WREADY,
  m_axi_in_10_WSTRB,
  m_axi_in_10_WVALID,
  m_axi_out_10_ARADDR,
  m_axi_out_10_ARBURST,
  m_axi_out_10_ARCACHE,
  m_axi_out_10_ARID,
  m_axi_out_10_ARLEN,
  m_axi_out_10_ARLOCK,
  m_axi_out_10_ARPROT,
  m_axi_out_10_ARQOS,
  m_axi_out_10_ARREADY,
  m_axi_out_10_ARSIZE,
  m_axi_out_10_ARVALID,
  m_axi_out_10_AWADDR,
  m_axi_out_10_AWBURST,
  m_axi_out_10_AWCACHE,
  m_axi_out_10_AWID,
  m_axi_out_10_AWLEN,
  m_axi_out_10_AWLOCK,
  m_axi_out_10_AWPROT,
  m_axi_out_10_AWQOS,
  m_axi_out_10_AWREADY,
  m_axi_out_10_AWSIZE,
  m_axi_out_10_AWVALID,
  m_axi_out_10_BID,
  m_axi_out_10_BREADY,
  m_axi_out_10_BRESP,
  m_axi_out_10_BVALID,
  m_axi_out_10_RDATA,
  m_axi_out_10_RID,
  m_axi_out_10_RLAST,
  m_axi_out_10_RREADY,
  m_axi_out_10_RRESP,
  m_axi_out_10_RVALID,
  m_axi_out_10_WDATA,
  m_axi_out_10_WLAST,
  m_axi_out_10_WREADY,
  m_axi_out_10_WSTRB,
  m_axi_out_10_WVALID,
  m_axi_in_11_ARADDR,
  m_axi_in_11_ARBURST,
  m_axi_in_11_ARCACHE,
  m_axi_in_11_ARID,
  m_axi_in_11_ARLEN,
  m_axi_in_11_ARLOCK,
  m_axi_in_11_ARPROT,
  m_axi_in_11_ARQOS,
  m_axi_in_11_ARREADY,
  m_axi_in_11_ARSIZE,
  m_axi_in_11_ARVALID,
  m_axi_in_11_AWADDR,
  m_axi_in_11_AWBURST,
  m_axi_in_11_AWCACHE,
  m_axi_in_11_AWID,
  m_axi_in_11_AWLEN,
  m_axi_in_11_AWLOCK,
  m_axi_in_11_AWPROT,
  m_axi_in_11_AWQOS,
  m_axi_in_11_AWREADY,
  m_axi_in_11_AWSIZE,
  m_axi_in_11_AWVALID,
  m_axi_in_11_BID,
  m_axi_in_11_BREADY,
  m_axi_in_11_BRESP,
  m_axi_in_11_BVALID,
  m_axi_in_11_RDATA,
  m_axi_in_11_RID,
  m_axi_in_11_RLAST,
  m_axi_in_11_RREADY,
  m_axi_in_11_RRESP,
  m_axi_in_11_RVALID,
  m_axi_in_11_WDATA,
  m_axi_in_11_WLAST,
  m_axi_in_11_WREADY,
  m_axi_in_11_WSTRB,
  m_axi_in_11_WVALID,
  m_axi_out_11_ARADDR,
  m_axi_out_11_ARBURST,
  m_axi_out_11_ARCACHE,
  m_axi_out_11_ARID,
  m_axi_out_11_ARLEN,
  m_axi_out_11_ARLOCK,
  m_axi_out_11_ARPROT,
  m_axi_out_11_ARQOS,
  m_axi_out_11_ARREADY,
  m_axi_out_11_ARSIZE,
  m_axi_out_11_ARVALID,
  m_axi_out_11_AWADDR,
  m_axi_out_11_AWBURST,
  m_axi_out_11_AWCACHE,
  m_axi_out_11_AWID,
  m_axi_out_11_AWLEN,
  m_axi_out_11_AWLOCK,
  m_axi_out_11_AWPROT,
  m_axi_out_11_AWQOS,
  m_axi_out_11_AWREADY,
  m_axi_out_11_AWSIZE,
  m_axi_out_11_AWVALID,
  m_axi_out_11_BID,
  m_axi_out_11_BREADY,
  m_axi_out_11_BRESP,
  m_axi_out_11_BVALID,
  m_axi_out_11_RDATA,
  m_axi_out_11_RID,
  m_axi_out_11_RLAST,
  m_axi_out_11_RREADY,
  m_axi_out_11_RRESP,
  m_axi_out_11_RVALID,
  m_axi_out_11_WDATA,
  m_axi_out_11_WLAST,
  m_axi_out_11_WREADY,
  m_axi_out_11_WSTRB,
  m_axi_out_11_WVALID,
  m_axi_in_12_ARADDR,
  m_axi_in_12_ARBURST,
  m_axi_in_12_ARCACHE,
  m_axi_in_12_ARID,
  m_axi_in_12_ARLEN,
  m_axi_in_12_ARLOCK,
  m_axi_in_12_ARPROT,
  m_axi_in_12_ARQOS,
  m_axi_in_12_ARREADY,
  m_axi_in_12_ARSIZE,
  m_axi_in_12_ARVALID,
  m_axi_in_12_AWADDR,
  m_axi_in_12_AWBURST,
  m_axi_in_12_AWCACHE,
  m_axi_in_12_AWID,
  m_axi_in_12_AWLEN,
  m_axi_in_12_AWLOCK,
  m_axi_in_12_AWPROT,
  m_axi_in_12_AWQOS,
  m_axi_in_12_AWREADY,
  m_axi_in_12_AWSIZE,
  m_axi_in_12_AWVALID,
  m_axi_in_12_BID,
  m_axi_in_12_BREADY,
  m_axi_in_12_BRESP,
  m_axi_in_12_BVALID,
  m_axi_in_12_RDATA,
  m_axi_in_12_RID,
  m_axi_in_12_RLAST,
  m_axi_in_12_RREADY,
  m_axi_in_12_RRESP,
  m_axi_in_12_RVALID,
  m_axi_in_12_WDATA,
  m_axi_in_12_WLAST,
  m_axi_in_12_WREADY,
  m_axi_in_12_WSTRB,
  m_axi_in_12_WVALID,
  m_axi_out_12_ARADDR,
  m_axi_out_12_ARBURST,
  m_axi_out_12_ARCACHE,
  m_axi_out_12_ARID,
  m_axi_out_12_ARLEN,
  m_axi_out_12_ARLOCK,
  m_axi_out_12_ARPROT,
  m_axi_out_12_ARQOS,
  m_axi_out_12_ARREADY,
  m_axi_out_12_ARSIZE,
  m_axi_out_12_ARVALID,
  m_axi_out_12_AWADDR,
  m_axi_out_12_AWBURST,
  m_axi_out_12_AWCACHE,
  m_axi_out_12_AWID,
  m_axi_out_12_AWLEN,
  m_axi_out_12_AWLOCK,
  m_axi_out_12_AWPROT,
  m_axi_out_12_AWQOS,
  m_axi_out_12_AWREADY,
  m_axi_out_12_AWSIZE,
  m_axi_out_12_AWVALID,
  m_axi_out_12_BID,
  m_axi_out_12_BREADY,
  m_axi_out_12_BRESP,
  m_axi_out_12_BVALID,
  m_axi_out_12_RDATA,
  m_axi_out_12_RID,
  m_axi_out_12_RLAST,
  m_axi_out_12_RREADY,
  m_axi_out_12_RRESP,
  m_axi_out_12_RVALID,
  m_axi_out_12_WDATA,
  m_axi_out_12_WLAST,
  m_axi_out_12_WREADY,
  m_axi_out_12_WSTRB,
  m_axi_out_12_WVALID,
  m_axi_in_13_ARADDR,
  m_axi_in_13_ARBURST,
  m_axi_in_13_ARCACHE,
  m_axi_in_13_ARID,
  m_axi_in_13_ARLEN,
  m_axi_in_13_ARLOCK,
  m_axi_in_13_ARPROT,
  m_axi_in_13_ARQOS,
  m_axi_in_13_ARREADY,
  m_axi_in_13_ARSIZE,
  m_axi_in_13_ARVALID,
  m_axi_in_13_AWADDR,
  m_axi_in_13_AWBURST,
  m_axi_in_13_AWCACHE,
  m_axi_in_13_AWID,
  m_axi_in_13_AWLEN,
  m_axi_in_13_AWLOCK,
  m_axi_in_13_AWPROT,
  m_axi_in_13_AWQOS,
  m_axi_in_13_AWREADY,
  m_axi_in_13_AWSIZE,
  m_axi_in_13_AWVALID,
  m_axi_in_13_BID,
  m_axi_in_13_BREADY,
  m_axi_in_13_BRESP,
  m_axi_in_13_BVALID,
  m_axi_in_13_RDATA,
  m_axi_in_13_RID,
  m_axi_in_13_RLAST,
  m_axi_in_13_RREADY,
  m_axi_in_13_RRESP,
  m_axi_in_13_RVALID,
  m_axi_in_13_WDATA,
  m_axi_in_13_WLAST,
  m_axi_in_13_WREADY,
  m_axi_in_13_WSTRB,
  m_axi_in_13_WVALID,
  m_axi_out_13_ARADDR,
  m_axi_out_13_ARBURST,
  m_axi_out_13_ARCACHE,
  m_axi_out_13_ARID,
  m_axi_out_13_ARLEN,
  m_axi_out_13_ARLOCK,
  m_axi_out_13_ARPROT,
  m_axi_out_13_ARQOS,
  m_axi_out_13_ARREADY,
  m_axi_out_13_ARSIZE,
  m_axi_out_13_ARVALID,
  m_axi_out_13_AWADDR,
  m_axi_out_13_AWBURST,
  m_axi_out_13_AWCACHE,
  m_axi_out_13_AWID,
  m_axi_out_13_AWLEN,
  m_axi_out_13_AWLOCK,
  m_axi_out_13_AWPROT,
  m_axi_out_13_AWQOS,
  m_axi_out_13_AWREADY,
  m_axi_out_13_AWSIZE,
  m_axi_out_13_AWVALID,
  m_axi_out_13_BID,
  m_axi_out_13_BREADY,
  m_axi_out_13_BRESP,
  m_axi_out_13_BVALID,
  m_axi_out_13_RDATA,
  m_axi_out_13_RID,
  m_axi_out_13_RLAST,
  m_axi_out_13_RREADY,
  m_axi_out_13_RRESP,
  m_axi_out_13_RVALID,
  m_axi_out_13_WDATA,
  m_axi_out_13_WLAST,
  m_axi_out_13_WREADY,
  m_axi_out_13_WSTRB,
  m_axi_out_13_WVALID,
  m_axi_in_14_ARADDR,
  m_axi_in_14_ARBURST,
  m_axi_in_14_ARCACHE,
  m_axi_in_14_ARID,
  m_axi_in_14_ARLEN,
  m_axi_in_14_ARLOCK,
  m_axi_in_14_ARPROT,
  m_axi_in_14_ARQOS,
  m_axi_in_14_ARREADY,
  m_axi_in_14_ARSIZE,
  m_axi_in_14_ARVALID,
  m_axi_in_14_AWADDR,
  m_axi_in_14_AWBURST,
  m_axi_in_14_AWCACHE,
  m_axi_in_14_AWID,
  m_axi_in_14_AWLEN,
  m_axi_in_14_AWLOCK,
  m_axi_in_14_AWPROT,
  m_axi_in_14_AWQOS,
  m_axi_in_14_AWREADY,
  m_axi_in_14_AWSIZE,
  m_axi_in_14_AWVALID,
  m_axi_in_14_BID,
  m_axi_in_14_BREADY,
  m_axi_in_14_BRESP,
  m_axi_in_14_BVALID,
  m_axi_in_14_RDATA,
  m_axi_in_14_RID,
  m_axi_in_14_RLAST,
  m_axi_in_14_RREADY,
  m_axi_in_14_RRESP,
  m_axi_in_14_RVALID,
  m_axi_in_14_WDATA,
  m_axi_in_14_WLAST,
  m_axi_in_14_WREADY,
  m_axi_in_14_WSTRB,
  m_axi_in_14_WVALID,
  m_axi_out_14_ARADDR,
  m_axi_out_14_ARBURST,
  m_axi_out_14_ARCACHE,
  m_axi_out_14_ARID,
  m_axi_out_14_ARLEN,
  m_axi_out_14_ARLOCK,
  m_axi_out_14_ARPROT,
  m_axi_out_14_ARQOS,
  m_axi_out_14_ARREADY,
  m_axi_out_14_ARSIZE,
  m_axi_out_14_ARVALID,
  m_axi_out_14_AWADDR,
  m_axi_out_14_AWBURST,
  m_axi_out_14_AWCACHE,
  m_axi_out_14_AWID,
  m_axi_out_14_AWLEN,
  m_axi_out_14_AWLOCK,
  m_axi_out_14_AWPROT,
  m_axi_out_14_AWQOS,
  m_axi_out_14_AWREADY,
  m_axi_out_14_AWSIZE,
  m_axi_out_14_AWVALID,
  m_axi_out_14_BID,
  m_axi_out_14_BREADY,
  m_axi_out_14_BRESP,
  m_axi_out_14_BVALID,
  m_axi_out_14_RDATA,
  m_axi_out_14_RID,
  m_axi_out_14_RLAST,
  m_axi_out_14_RREADY,
  m_axi_out_14_RRESP,
  m_axi_out_14_RVALID,
  m_axi_out_14_WDATA,
  m_axi_out_14_WLAST,
  m_axi_out_14_WREADY,
  m_axi_out_14_WSTRB,
  m_axi_out_14_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 9;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  (* RS_HS = "s_axi_control_AW.valid" *)input s_axi_control_AWVALID;
  (* RS_HS = "s_axi_control_AW.ready" *)output s_axi_control_AWREADY;
  (* RS_HS = "s_axi_control_AW.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  (* RS_HS = "s_axi_control_W.valid" *)input s_axi_control_WVALID;
  (* RS_HS = "s_axi_control_W.ready" *)output s_axi_control_WREADY;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  (* RS_HS = "s_axi_control_AR.valid" *)input s_axi_control_ARVALID;
  (* RS_HS = "s_axi_control_AR.ready" *)output s_axi_control_ARREADY;
  (* RS_HS = "s_axi_control_AR.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  (* RS_HS = "s_axi_control_R.valid" *)output s_axi_control_RVALID;
  (* RS_HS = "s_axi_control_R.ready" *)input s_axi_control_RREADY;
  (* RS_HS = "s_axi_control_R.data" *)output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  (* RS_HS = "s_axi_control_R.data" *)output [1:0] s_axi_control_RRESP;
  (* RS_HS = "s_axi_control_B.valid" *)output s_axi_control_BVALID;
  (* RS_HS = "s_axi_control_B.ready" *)input s_axi_control_BREADY;
  (* RS_HS = "s_axi_control_B.data" *)output [1:0] s_axi_control_BRESP;
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_FF = "interrupt" *)output interrupt;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [63:0] m_axi_in_0_ARADDR;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [1:0] m_axi_in_0_ARBURST;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [3:0] m_axi_in_0_ARCACHE;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [0:0] m_axi_in_0_ARID;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [7:0] m_axi_in_0_ARLEN;
  (* RS_HS = "m_axi_in_0_AR.data" *)output m_axi_in_0_ARLOCK;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [2:0] m_axi_in_0_ARPROT;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [3:0] m_axi_in_0_ARQOS;
  (* RS_HS = "m_axi_in_0_AR.ready" *)input m_axi_in_0_ARREADY;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [2:0] m_axi_in_0_ARSIZE;
  (* RS_HS = "m_axi_in_0_AR.valid" *)output m_axi_in_0_ARVALID;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [63:0] m_axi_in_0_AWADDR;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [1:0] m_axi_in_0_AWBURST;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [3:0] m_axi_in_0_AWCACHE;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [0:0] m_axi_in_0_AWID;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [7:0] m_axi_in_0_AWLEN;
  (* RS_HS = "m_axi_in_0_AW.data" *)output m_axi_in_0_AWLOCK;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [2:0] m_axi_in_0_AWPROT;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [3:0] m_axi_in_0_AWQOS;
  (* RS_HS = "m_axi_in_0_AW.ready" *)input m_axi_in_0_AWREADY;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [2:0] m_axi_in_0_AWSIZE;
  (* RS_HS = "m_axi_in_0_AW.valid" *)output m_axi_in_0_AWVALID;
  (* RS_HS = "m_axi_in_0_B.data" *)input [0:0] m_axi_in_0_BID;
  (* RS_HS = "m_axi_in_0_B.ready" *)output m_axi_in_0_BREADY;
  (* RS_HS = "m_axi_in_0_B.data" *)input [1:0] m_axi_in_0_BRESP;
  (* RS_HS = "m_axi_in_0_B.valid" *)input m_axi_in_0_BVALID;
  (* RS_HS = "m_axi_in_0_R.data" *)input [511:0] m_axi_in_0_RDATA;
  (* RS_HS = "m_axi_in_0_R.data" *)input [0:0] m_axi_in_0_RID;
  (* RS_HS = "m_axi_in_0_R.data" *)input m_axi_in_0_RLAST;
  (* RS_HS = "m_axi_in_0_R.ready" *)output m_axi_in_0_RREADY;
  (* RS_HS = "m_axi_in_0_R.data" *)input [1:0] m_axi_in_0_RRESP;
  (* RS_HS = "m_axi_in_0_R.valid" *)input m_axi_in_0_RVALID;
  (* RS_HS = "m_axi_in_0_W.data" *)output [511:0] m_axi_in_0_WDATA;
  (* RS_HS = "m_axi_in_0_W.data" *)output m_axi_in_0_WLAST;
  (* RS_HS = "m_axi_in_0_W.ready" *)input m_axi_in_0_WREADY;
  (* RS_HS = "m_axi_in_0_W.data" *)output [63:0] m_axi_in_0_WSTRB;
  (* RS_HS = "m_axi_in_0_W.valid" *)output m_axi_in_0_WVALID;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [63:0] m_axi_out_0_ARADDR;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [1:0] m_axi_out_0_ARBURST;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [3:0] m_axi_out_0_ARCACHE;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [0:0] m_axi_out_0_ARID;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [7:0] m_axi_out_0_ARLEN;
  (* RS_HS = "m_axi_out_0_AR.data" *)output m_axi_out_0_ARLOCK;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [2:0] m_axi_out_0_ARPROT;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [3:0] m_axi_out_0_ARQOS;
  (* RS_HS = "m_axi_out_0_AR.ready" *)input m_axi_out_0_ARREADY;
  (* RS_HS = "m_axi_out_0_AR.data" *)output [2:0] m_axi_out_0_ARSIZE;
  (* RS_HS = "m_axi_out_0_AR.valid" *)output m_axi_out_0_ARVALID;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [63:0] m_axi_out_0_AWADDR;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [1:0] m_axi_out_0_AWBURST;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [3:0] m_axi_out_0_AWCACHE;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [0:0] m_axi_out_0_AWID;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [7:0] m_axi_out_0_AWLEN;
  (* RS_HS = "m_axi_out_0_AW.data" *)output m_axi_out_0_AWLOCK;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [2:0] m_axi_out_0_AWPROT;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [3:0] m_axi_out_0_AWQOS;
  (* RS_HS = "m_axi_out_0_AW.ready" *)input m_axi_out_0_AWREADY;
  (* RS_HS = "m_axi_out_0_AW.data" *)output [2:0] m_axi_out_0_AWSIZE;
  (* RS_HS = "m_axi_out_0_AW.valid" *)output m_axi_out_0_AWVALID;
  (* RS_HS = "m_axi_out_0_B.data" *)input [0:0] m_axi_out_0_BID;
  (* RS_HS = "m_axi_out_0_B.ready" *)output m_axi_out_0_BREADY;
  (* RS_HS = "m_axi_out_0_B.data" *)input [1:0] m_axi_out_0_BRESP;
  (* RS_HS = "m_axi_out_0_B.valid" *)input m_axi_out_0_BVALID;
  (* RS_HS = "m_axi_out_0_R.data" *)input [511:0] m_axi_out_0_RDATA;
  (* RS_HS = "m_axi_out_0_R.data" *)input [0:0] m_axi_out_0_RID;
  (* RS_HS = "m_axi_out_0_R.data" *)input m_axi_out_0_RLAST;
  (* RS_HS = "m_axi_out_0_R.ready" *)output m_axi_out_0_RREADY;
  (* RS_HS = "m_axi_out_0_R.data" *)input [1:0] m_axi_out_0_RRESP;
  (* RS_HS = "m_axi_out_0_R.valid" *)input m_axi_out_0_RVALID;
  (* RS_HS = "m_axi_out_0_W.data" *)output [511:0] m_axi_out_0_WDATA;
  (* RS_HS = "m_axi_out_0_W.data" *)output m_axi_out_0_WLAST;
  (* RS_HS = "m_axi_out_0_W.ready" *)input m_axi_out_0_WREADY;
  (* RS_HS = "m_axi_out_0_W.data" *)output [63:0] m_axi_out_0_WSTRB;
  (* RS_HS = "m_axi_out_0_W.valid" *)output m_axi_out_0_WVALID;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [63:0] m_axi_in_1_ARADDR;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [1:0] m_axi_in_1_ARBURST;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [3:0] m_axi_in_1_ARCACHE;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [0:0] m_axi_in_1_ARID;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [7:0] m_axi_in_1_ARLEN;
  (* RS_HS = "m_axi_in_1_AR.data" *)output m_axi_in_1_ARLOCK;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [2:0] m_axi_in_1_ARPROT;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [3:0] m_axi_in_1_ARQOS;
  (* RS_HS = "m_axi_in_1_AR.ready" *)input m_axi_in_1_ARREADY;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [2:0] m_axi_in_1_ARSIZE;
  (* RS_HS = "m_axi_in_1_AR.valid" *)output m_axi_in_1_ARVALID;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [63:0] m_axi_in_1_AWADDR;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [1:0] m_axi_in_1_AWBURST;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [3:0] m_axi_in_1_AWCACHE;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [0:0] m_axi_in_1_AWID;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [7:0] m_axi_in_1_AWLEN;
  (* RS_HS = "m_axi_in_1_AW.data" *)output m_axi_in_1_AWLOCK;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [2:0] m_axi_in_1_AWPROT;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [3:0] m_axi_in_1_AWQOS;
  (* RS_HS = "m_axi_in_1_AW.ready" *)input m_axi_in_1_AWREADY;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [2:0] m_axi_in_1_AWSIZE;
  (* RS_HS = "m_axi_in_1_AW.valid" *)output m_axi_in_1_AWVALID;
  (* RS_HS = "m_axi_in_1_B.data" *)input [0:0] m_axi_in_1_BID;
  (* RS_HS = "m_axi_in_1_B.ready" *)output m_axi_in_1_BREADY;
  (* RS_HS = "m_axi_in_1_B.data" *)input [1:0] m_axi_in_1_BRESP;
  (* RS_HS = "m_axi_in_1_B.valid" *)input m_axi_in_1_BVALID;
  (* RS_HS = "m_axi_in_1_R.data" *)input [511:0] m_axi_in_1_RDATA;
  (* RS_HS = "m_axi_in_1_R.data" *)input [0:0] m_axi_in_1_RID;
  (* RS_HS = "m_axi_in_1_R.data" *)input m_axi_in_1_RLAST;
  (* RS_HS = "m_axi_in_1_R.ready" *)output m_axi_in_1_RREADY;
  (* RS_HS = "m_axi_in_1_R.data" *)input [1:0] m_axi_in_1_RRESP;
  (* RS_HS = "m_axi_in_1_R.valid" *)input m_axi_in_1_RVALID;
  (* RS_HS = "m_axi_in_1_W.data" *)output [511:0] m_axi_in_1_WDATA;
  (* RS_HS = "m_axi_in_1_W.data" *)output m_axi_in_1_WLAST;
  (* RS_HS = "m_axi_in_1_W.ready" *)input m_axi_in_1_WREADY;
  (* RS_HS = "m_axi_in_1_W.data" *)output [63:0] m_axi_in_1_WSTRB;
  (* RS_HS = "m_axi_in_1_W.valid" *)output m_axi_in_1_WVALID;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [63:0] m_axi_out_1_ARADDR;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [1:0] m_axi_out_1_ARBURST;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [3:0] m_axi_out_1_ARCACHE;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [0:0] m_axi_out_1_ARID;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [7:0] m_axi_out_1_ARLEN;
  (* RS_HS = "m_axi_out_1_AR.data" *)output m_axi_out_1_ARLOCK;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [2:0] m_axi_out_1_ARPROT;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [3:0] m_axi_out_1_ARQOS;
  (* RS_HS = "m_axi_out_1_AR.ready" *)input m_axi_out_1_ARREADY;
  (* RS_HS = "m_axi_out_1_AR.data" *)output [2:0] m_axi_out_1_ARSIZE;
  (* RS_HS = "m_axi_out_1_AR.valid" *)output m_axi_out_1_ARVALID;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [63:0] m_axi_out_1_AWADDR;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [1:0] m_axi_out_1_AWBURST;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [3:0] m_axi_out_1_AWCACHE;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [0:0] m_axi_out_1_AWID;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [7:0] m_axi_out_1_AWLEN;
  (* RS_HS = "m_axi_out_1_AW.data" *)output m_axi_out_1_AWLOCK;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [2:0] m_axi_out_1_AWPROT;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [3:0] m_axi_out_1_AWQOS;
  (* RS_HS = "m_axi_out_1_AW.ready" *)input m_axi_out_1_AWREADY;
  (* RS_HS = "m_axi_out_1_AW.data" *)output [2:0] m_axi_out_1_AWSIZE;
  (* RS_HS = "m_axi_out_1_AW.valid" *)output m_axi_out_1_AWVALID;
  (* RS_HS = "m_axi_out_1_B.data" *)input [0:0] m_axi_out_1_BID;
  (* RS_HS = "m_axi_out_1_B.ready" *)output m_axi_out_1_BREADY;
  (* RS_HS = "m_axi_out_1_B.data" *)input [1:0] m_axi_out_1_BRESP;
  (* RS_HS = "m_axi_out_1_B.valid" *)input m_axi_out_1_BVALID;
  (* RS_HS = "m_axi_out_1_R.data" *)input [511:0] m_axi_out_1_RDATA;
  (* RS_HS = "m_axi_out_1_R.data" *)input [0:0] m_axi_out_1_RID;
  (* RS_HS = "m_axi_out_1_R.data" *)input m_axi_out_1_RLAST;
  (* RS_HS = "m_axi_out_1_R.ready" *)output m_axi_out_1_RREADY;
  (* RS_HS = "m_axi_out_1_R.data" *)input [1:0] m_axi_out_1_RRESP;
  (* RS_HS = "m_axi_out_1_R.valid" *)input m_axi_out_1_RVALID;
  (* RS_HS = "m_axi_out_1_W.data" *)output [511:0] m_axi_out_1_WDATA;
  (* RS_HS = "m_axi_out_1_W.data" *)output m_axi_out_1_WLAST;
  (* RS_HS = "m_axi_out_1_W.ready" *)input m_axi_out_1_WREADY;
  (* RS_HS = "m_axi_out_1_W.data" *)output [63:0] m_axi_out_1_WSTRB;
  (* RS_HS = "m_axi_out_1_W.valid" *)output m_axi_out_1_WVALID;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [63:0] m_axi_in_2_ARADDR;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [1:0] m_axi_in_2_ARBURST;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [3:0] m_axi_in_2_ARCACHE;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [0:0] m_axi_in_2_ARID;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [7:0] m_axi_in_2_ARLEN;
  (* RS_HS = "m_axi_in_2_AR.data" *)output m_axi_in_2_ARLOCK;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [2:0] m_axi_in_2_ARPROT;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [3:0] m_axi_in_2_ARQOS;
  (* RS_HS = "m_axi_in_2_AR.ready" *)input m_axi_in_2_ARREADY;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [2:0] m_axi_in_2_ARSIZE;
  (* RS_HS = "m_axi_in_2_AR.valid" *)output m_axi_in_2_ARVALID;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [63:0] m_axi_in_2_AWADDR;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [1:0] m_axi_in_2_AWBURST;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [3:0] m_axi_in_2_AWCACHE;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [0:0] m_axi_in_2_AWID;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [7:0] m_axi_in_2_AWLEN;
  (* RS_HS = "m_axi_in_2_AW.data" *)output m_axi_in_2_AWLOCK;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [2:0] m_axi_in_2_AWPROT;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [3:0] m_axi_in_2_AWQOS;
  (* RS_HS = "m_axi_in_2_AW.ready" *)input m_axi_in_2_AWREADY;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [2:0] m_axi_in_2_AWSIZE;
  (* RS_HS = "m_axi_in_2_AW.valid" *)output m_axi_in_2_AWVALID;
  (* RS_HS = "m_axi_in_2_B.data" *)input [0:0] m_axi_in_2_BID;
  (* RS_HS = "m_axi_in_2_B.ready" *)output m_axi_in_2_BREADY;
  (* RS_HS = "m_axi_in_2_B.data" *)input [1:0] m_axi_in_2_BRESP;
  (* RS_HS = "m_axi_in_2_B.valid" *)input m_axi_in_2_BVALID;
  (* RS_HS = "m_axi_in_2_R.data" *)input [511:0] m_axi_in_2_RDATA;
  (* RS_HS = "m_axi_in_2_R.data" *)input [0:0] m_axi_in_2_RID;
  (* RS_HS = "m_axi_in_2_R.data" *)input m_axi_in_2_RLAST;
  (* RS_HS = "m_axi_in_2_R.ready" *)output m_axi_in_2_RREADY;
  (* RS_HS = "m_axi_in_2_R.data" *)input [1:0] m_axi_in_2_RRESP;
  (* RS_HS = "m_axi_in_2_R.valid" *)input m_axi_in_2_RVALID;
  (* RS_HS = "m_axi_in_2_W.data" *)output [511:0] m_axi_in_2_WDATA;
  (* RS_HS = "m_axi_in_2_W.data" *)output m_axi_in_2_WLAST;
  (* RS_HS = "m_axi_in_2_W.ready" *)input m_axi_in_2_WREADY;
  (* RS_HS = "m_axi_in_2_W.data" *)output [63:0] m_axi_in_2_WSTRB;
  (* RS_HS = "m_axi_in_2_W.valid" *)output m_axi_in_2_WVALID;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [63:0] m_axi_out_2_ARADDR;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [1:0] m_axi_out_2_ARBURST;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [3:0] m_axi_out_2_ARCACHE;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [0:0] m_axi_out_2_ARID;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [7:0] m_axi_out_2_ARLEN;
  (* RS_HS = "m_axi_out_2_AR.data" *)output m_axi_out_2_ARLOCK;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [2:0] m_axi_out_2_ARPROT;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [3:0] m_axi_out_2_ARQOS;
  (* RS_HS = "m_axi_out_2_AR.ready" *)input m_axi_out_2_ARREADY;
  (* RS_HS = "m_axi_out_2_AR.data" *)output [2:0] m_axi_out_2_ARSIZE;
  (* RS_HS = "m_axi_out_2_AR.valid" *)output m_axi_out_2_ARVALID;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [63:0] m_axi_out_2_AWADDR;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [1:0] m_axi_out_2_AWBURST;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [3:0] m_axi_out_2_AWCACHE;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [0:0] m_axi_out_2_AWID;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [7:0] m_axi_out_2_AWLEN;
  (* RS_HS = "m_axi_out_2_AW.data" *)output m_axi_out_2_AWLOCK;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [2:0] m_axi_out_2_AWPROT;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [3:0] m_axi_out_2_AWQOS;
  (* RS_HS = "m_axi_out_2_AW.ready" *)input m_axi_out_2_AWREADY;
  (* RS_HS = "m_axi_out_2_AW.data" *)output [2:0] m_axi_out_2_AWSIZE;
  (* RS_HS = "m_axi_out_2_AW.valid" *)output m_axi_out_2_AWVALID;
  (* RS_HS = "m_axi_out_2_B.data" *)input [0:0] m_axi_out_2_BID;
  (* RS_HS = "m_axi_out_2_B.ready" *)output m_axi_out_2_BREADY;
  (* RS_HS = "m_axi_out_2_B.data" *)input [1:0] m_axi_out_2_BRESP;
  (* RS_HS = "m_axi_out_2_B.valid" *)input m_axi_out_2_BVALID;
  (* RS_HS = "m_axi_out_2_R.data" *)input [511:0] m_axi_out_2_RDATA;
  (* RS_HS = "m_axi_out_2_R.data" *)input [0:0] m_axi_out_2_RID;
  (* RS_HS = "m_axi_out_2_R.data" *)input m_axi_out_2_RLAST;
  (* RS_HS = "m_axi_out_2_R.ready" *)output m_axi_out_2_RREADY;
  (* RS_HS = "m_axi_out_2_R.data" *)input [1:0] m_axi_out_2_RRESP;
  (* RS_HS = "m_axi_out_2_R.valid" *)input m_axi_out_2_RVALID;
  (* RS_HS = "m_axi_out_2_W.data" *)output [511:0] m_axi_out_2_WDATA;
  (* RS_HS = "m_axi_out_2_W.data" *)output m_axi_out_2_WLAST;
  (* RS_HS = "m_axi_out_2_W.ready" *)input m_axi_out_2_WREADY;
  (* RS_HS = "m_axi_out_2_W.data" *)output [63:0] m_axi_out_2_WSTRB;
  (* RS_HS = "m_axi_out_2_W.valid" *)output m_axi_out_2_WVALID;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [63:0] m_axi_in_3_ARADDR;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [1:0] m_axi_in_3_ARBURST;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [3:0] m_axi_in_3_ARCACHE;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [0:0] m_axi_in_3_ARID;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [7:0] m_axi_in_3_ARLEN;
  (* RS_HS = "m_axi_in_3_AR.data" *)output m_axi_in_3_ARLOCK;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [2:0] m_axi_in_3_ARPROT;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [3:0] m_axi_in_3_ARQOS;
  (* RS_HS = "m_axi_in_3_AR.ready" *)input m_axi_in_3_ARREADY;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [2:0] m_axi_in_3_ARSIZE;
  (* RS_HS = "m_axi_in_3_AR.valid" *)output m_axi_in_3_ARVALID;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [63:0] m_axi_in_3_AWADDR;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [1:0] m_axi_in_3_AWBURST;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [3:0] m_axi_in_3_AWCACHE;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [0:0] m_axi_in_3_AWID;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [7:0] m_axi_in_3_AWLEN;
  (* RS_HS = "m_axi_in_3_AW.data" *)output m_axi_in_3_AWLOCK;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [2:0] m_axi_in_3_AWPROT;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [3:0] m_axi_in_3_AWQOS;
  (* RS_HS = "m_axi_in_3_AW.ready" *)input m_axi_in_3_AWREADY;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [2:0] m_axi_in_3_AWSIZE;
  (* RS_HS = "m_axi_in_3_AW.valid" *)output m_axi_in_3_AWVALID;
  (* RS_HS = "m_axi_in_3_B.data" *)input [0:0] m_axi_in_3_BID;
  (* RS_HS = "m_axi_in_3_B.ready" *)output m_axi_in_3_BREADY;
  (* RS_HS = "m_axi_in_3_B.data" *)input [1:0] m_axi_in_3_BRESP;
  (* RS_HS = "m_axi_in_3_B.valid" *)input m_axi_in_3_BVALID;
  (* RS_HS = "m_axi_in_3_R.data" *)input [511:0] m_axi_in_3_RDATA;
  (* RS_HS = "m_axi_in_3_R.data" *)input [0:0] m_axi_in_3_RID;
  (* RS_HS = "m_axi_in_3_R.data" *)input m_axi_in_3_RLAST;
  (* RS_HS = "m_axi_in_3_R.ready" *)output m_axi_in_3_RREADY;
  (* RS_HS = "m_axi_in_3_R.data" *)input [1:0] m_axi_in_3_RRESP;
  (* RS_HS = "m_axi_in_3_R.valid" *)input m_axi_in_3_RVALID;
  (* RS_HS = "m_axi_in_3_W.data" *)output [511:0] m_axi_in_3_WDATA;
  (* RS_HS = "m_axi_in_3_W.data" *)output m_axi_in_3_WLAST;
  (* RS_HS = "m_axi_in_3_W.ready" *)input m_axi_in_3_WREADY;
  (* RS_HS = "m_axi_in_3_W.data" *)output [63:0] m_axi_in_3_WSTRB;
  (* RS_HS = "m_axi_in_3_W.valid" *)output m_axi_in_3_WVALID;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [63:0] m_axi_out_3_ARADDR;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [1:0] m_axi_out_3_ARBURST;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [3:0] m_axi_out_3_ARCACHE;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [0:0] m_axi_out_3_ARID;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [7:0] m_axi_out_3_ARLEN;
  (* RS_HS = "m_axi_out_3_AR.data" *)output m_axi_out_3_ARLOCK;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [2:0] m_axi_out_3_ARPROT;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [3:0] m_axi_out_3_ARQOS;
  (* RS_HS = "m_axi_out_3_AR.ready" *)input m_axi_out_3_ARREADY;
  (* RS_HS = "m_axi_out_3_AR.data" *)output [2:0] m_axi_out_3_ARSIZE;
  (* RS_HS = "m_axi_out_3_AR.valid" *)output m_axi_out_3_ARVALID;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [63:0] m_axi_out_3_AWADDR;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [1:0] m_axi_out_3_AWBURST;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [3:0] m_axi_out_3_AWCACHE;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [0:0] m_axi_out_3_AWID;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [7:0] m_axi_out_3_AWLEN;
  (* RS_HS = "m_axi_out_3_AW.data" *)output m_axi_out_3_AWLOCK;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [2:0] m_axi_out_3_AWPROT;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [3:0] m_axi_out_3_AWQOS;
  (* RS_HS = "m_axi_out_3_AW.ready" *)input m_axi_out_3_AWREADY;
  (* RS_HS = "m_axi_out_3_AW.data" *)output [2:0] m_axi_out_3_AWSIZE;
  (* RS_HS = "m_axi_out_3_AW.valid" *)output m_axi_out_3_AWVALID;
  (* RS_HS = "m_axi_out_3_B.data" *)input [0:0] m_axi_out_3_BID;
  (* RS_HS = "m_axi_out_3_B.ready" *)output m_axi_out_3_BREADY;
  (* RS_HS = "m_axi_out_3_B.data" *)input [1:0] m_axi_out_3_BRESP;
  (* RS_HS = "m_axi_out_3_B.valid" *)input m_axi_out_3_BVALID;
  (* RS_HS = "m_axi_out_3_R.data" *)input [511:0] m_axi_out_3_RDATA;
  (* RS_HS = "m_axi_out_3_R.data" *)input [0:0] m_axi_out_3_RID;
  (* RS_HS = "m_axi_out_3_R.data" *)input m_axi_out_3_RLAST;
  (* RS_HS = "m_axi_out_3_R.ready" *)output m_axi_out_3_RREADY;
  (* RS_HS = "m_axi_out_3_R.data" *)input [1:0] m_axi_out_3_RRESP;
  (* RS_HS = "m_axi_out_3_R.valid" *)input m_axi_out_3_RVALID;
  (* RS_HS = "m_axi_out_3_W.data" *)output [511:0] m_axi_out_3_WDATA;
  (* RS_HS = "m_axi_out_3_W.data" *)output m_axi_out_3_WLAST;
  (* RS_HS = "m_axi_out_3_W.ready" *)input m_axi_out_3_WREADY;
  (* RS_HS = "m_axi_out_3_W.data" *)output [63:0] m_axi_out_3_WSTRB;
  (* RS_HS = "m_axi_out_3_W.valid" *)output m_axi_out_3_WVALID;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [63:0] m_axi_in_4_ARADDR;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [1:0] m_axi_in_4_ARBURST;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [3:0] m_axi_in_4_ARCACHE;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [0:0] m_axi_in_4_ARID;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [7:0] m_axi_in_4_ARLEN;
  (* RS_HS = "m_axi_in_4_AR.data" *)output m_axi_in_4_ARLOCK;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [2:0] m_axi_in_4_ARPROT;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [3:0] m_axi_in_4_ARQOS;
  (* RS_HS = "m_axi_in_4_AR.ready" *)input m_axi_in_4_ARREADY;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [2:0] m_axi_in_4_ARSIZE;
  (* RS_HS = "m_axi_in_4_AR.valid" *)output m_axi_in_4_ARVALID;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [63:0] m_axi_in_4_AWADDR;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [1:0] m_axi_in_4_AWBURST;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [3:0] m_axi_in_4_AWCACHE;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [0:0] m_axi_in_4_AWID;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [7:0] m_axi_in_4_AWLEN;
  (* RS_HS = "m_axi_in_4_AW.data" *)output m_axi_in_4_AWLOCK;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [2:0] m_axi_in_4_AWPROT;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [3:0] m_axi_in_4_AWQOS;
  (* RS_HS = "m_axi_in_4_AW.ready" *)input m_axi_in_4_AWREADY;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [2:0] m_axi_in_4_AWSIZE;
  (* RS_HS = "m_axi_in_4_AW.valid" *)output m_axi_in_4_AWVALID;
  (* RS_HS = "m_axi_in_4_B.data" *)input [0:0] m_axi_in_4_BID;
  (* RS_HS = "m_axi_in_4_B.ready" *)output m_axi_in_4_BREADY;
  (* RS_HS = "m_axi_in_4_B.data" *)input [1:0] m_axi_in_4_BRESP;
  (* RS_HS = "m_axi_in_4_B.valid" *)input m_axi_in_4_BVALID;
  (* RS_HS = "m_axi_in_4_R.data" *)input [511:0] m_axi_in_4_RDATA;
  (* RS_HS = "m_axi_in_4_R.data" *)input [0:0] m_axi_in_4_RID;
  (* RS_HS = "m_axi_in_4_R.data" *)input m_axi_in_4_RLAST;
  (* RS_HS = "m_axi_in_4_R.ready" *)output m_axi_in_4_RREADY;
  (* RS_HS = "m_axi_in_4_R.data" *)input [1:0] m_axi_in_4_RRESP;
  (* RS_HS = "m_axi_in_4_R.valid" *)input m_axi_in_4_RVALID;
  (* RS_HS = "m_axi_in_4_W.data" *)output [511:0] m_axi_in_4_WDATA;
  (* RS_HS = "m_axi_in_4_W.data" *)output m_axi_in_4_WLAST;
  (* RS_HS = "m_axi_in_4_W.ready" *)input m_axi_in_4_WREADY;
  (* RS_HS = "m_axi_in_4_W.data" *)output [63:0] m_axi_in_4_WSTRB;
  (* RS_HS = "m_axi_in_4_W.valid" *)output m_axi_in_4_WVALID;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [63:0] m_axi_out_4_ARADDR;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [1:0] m_axi_out_4_ARBURST;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [3:0] m_axi_out_4_ARCACHE;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [0:0] m_axi_out_4_ARID;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [7:0] m_axi_out_4_ARLEN;
  (* RS_HS = "m_axi_out_4_AR.data" *)output m_axi_out_4_ARLOCK;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [2:0] m_axi_out_4_ARPROT;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [3:0] m_axi_out_4_ARQOS;
  (* RS_HS = "m_axi_out_4_AR.ready" *)input m_axi_out_4_ARREADY;
  (* RS_HS = "m_axi_out_4_AR.data" *)output [2:0] m_axi_out_4_ARSIZE;
  (* RS_HS = "m_axi_out_4_AR.valid" *)output m_axi_out_4_ARVALID;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [63:0] m_axi_out_4_AWADDR;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [1:0] m_axi_out_4_AWBURST;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [3:0] m_axi_out_4_AWCACHE;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [0:0] m_axi_out_4_AWID;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [7:0] m_axi_out_4_AWLEN;
  (* RS_HS = "m_axi_out_4_AW.data" *)output m_axi_out_4_AWLOCK;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [2:0] m_axi_out_4_AWPROT;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [3:0] m_axi_out_4_AWQOS;
  (* RS_HS = "m_axi_out_4_AW.ready" *)input m_axi_out_4_AWREADY;
  (* RS_HS = "m_axi_out_4_AW.data" *)output [2:0] m_axi_out_4_AWSIZE;
  (* RS_HS = "m_axi_out_4_AW.valid" *)output m_axi_out_4_AWVALID;
  (* RS_HS = "m_axi_out_4_B.data" *)input [0:0] m_axi_out_4_BID;
  (* RS_HS = "m_axi_out_4_B.ready" *)output m_axi_out_4_BREADY;
  (* RS_HS = "m_axi_out_4_B.data" *)input [1:0] m_axi_out_4_BRESP;
  (* RS_HS = "m_axi_out_4_B.valid" *)input m_axi_out_4_BVALID;
  (* RS_HS = "m_axi_out_4_R.data" *)input [511:0] m_axi_out_4_RDATA;
  (* RS_HS = "m_axi_out_4_R.data" *)input [0:0] m_axi_out_4_RID;
  (* RS_HS = "m_axi_out_4_R.data" *)input m_axi_out_4_RLAST;
  (* RS_HS = "m_axi_out_4_R.ready" *)output m_axi_out_4_RREADY;
  (* RS_HS = "m_axi_out_4_R.data" *)input [1:0] m_axi_out_4_RRESP;
  (* RS_HS = "m_axi_out_4_R.valid" *)input m_axi_out_4_RVALID;
  (* RS_HS = "m_axi_out_4_W.data" *)output [511:0] m_axi_out_4_WDATA;
  (* RS_HS = "m_axi_out_4_W.data" *)output m_axi_out_4_WLAST;
  (* RS_HS = "m_axi_out_4_W.ready" *)input m_axi_out_4_WREADY;
  (* RS_HS = "m_axi_out_4_W.data" *)output [63:0] m_axi_out_4_WSTRB;
  (* RS_HS = "m_axi_out_4_W.valid" *)output m_axi_out_4_WVALID;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [63:0] m_axi_in_5_ARADDR;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [1:0] m_axi_in_5_ARBURST;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [3:0] m_axi_in_5_ARCACHE;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [0:0] m_axi_in_5_ARID;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [7:0] m_axi_in_5_ARLEN;
  (* RS_HS = "m_axi_in_5_AR.data" *)output m_axi_in_5_ARLOCK;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [2:0] m_axi_in_5_ARPROT;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [3:0] m_axi_in_5_ARQOS;
  (* RS_HS = "m_axi_in_5_AR.ready" *)input m_axi_in_5_ARREADY;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [2:0] m_axi_in_5_ARSIZE;
  (* RS_HS = "m_axi_in_5_AR.valid" *)output m_axi_in_5_ARVALID;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [63:0] m_axi_in_5_AWADDR;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [1:0] m_axi_in_5_AWBURST;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [3:0] m_axi_in_5_AWCACHE;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [0:0] m_axi_in_5_AWID;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [7:0] m_axi_in_5_AWLEN;
  (* RS_HS = "m_axi_in_5_AW.data" *)output m_axi_in_5_AWLOCK;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [2:0] m_axi_in_5_AWPROT;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [3:0] m_axi_in_5_AWQOS;
  (* RS_HS = "m_axi_in_5_AW.ready" *)input m_axi_in_5_AWREADY;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [2:0] m_axi_in_5_AWSIZE;
  (* RS_HS = "m_axi_in_5_AW.valid" *)output m_axi_in_5_AWVALID;
  (* RS_HS = "m_axi_in_5_B.data" *)input [0:0] m_axi_in_5_BID;
  (* RS_HS = "m_axi_in_5_B.ready" *)output m_axi_in_5_BREADY;
  (* RS_HS = "m_axi_in_5_B.data" *)input [1:0] m_axi_in_5_BRESP;
  (* RS_HS = "m_axi_in_5_B.valid" *)input m_axi_in_5_BVALID;
  (* RS_HS = "m_axi_in_5_R.data" *)input [511:0] m_axi_in_5_RDATA;
  (* RS_HS = "m_axi_in_5_R.data" *)input [0:0] m_axi_in_5_RID;
  (* RS_HS = "m_axi_in_5_R.data" *)input m_axi_in_5_RLAST;
  (* RS_HS = "m_axi_in_5_R.ready" *)output m_axi_in_5_RREADY;
  (* RS_HS = "m_axi_in_5_R.data" *)input [1:0] m_axi_in_5_RRESP;
  (* RS_HS = "m_axi_in_5_R.valid" *)input m_axi_in_5_RVALID;
  (* RS_HS = "m_axi_in_5_W.data" *)output [511:0] m_axi_in_5_WDATA;
  (* RS_HS = "m_axi_in_5_W.data" *)output m_axi_in_5_WLAST;
  (* RS_HS = "m_axi_in_5_W.ready" *)input m_axi_in_5_WREADY;
  (* RS_HS = "m_axi_in_5_W.data" *)output [63:0] m_axi_in_5_WSTRB;
  (* RS_HS = "m_axi_in_5_W.valid" *)output m_axi_in_5_WVALID;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [63:0] m_axi_out_5_ARADDR;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [1:0] m_axi_out_5_ARBURST;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [3:0] m_axi_out_5_ARCACHE;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [0:0] m_axi_out_5_ARID;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [7:0] m_axi_out_5_ARLEN;
  (* RS_HS = "m_axi_out_5_AR.data" *)output m_axi_out_5_ARLOCK;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [2:0] m_axi_out_5_ARPROT;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [3:0] m_axi_out_5_ARQOS;
  (* RS_HS = "m_axi_out_5_AR.ready" *)input m_axi_out_5_ARREADY;
  (* RS_HS = "m_axi_out_5_AR.data" *)output [2:0] m_axi_out_5_ARSIZE;
  (* RS_HS = "m_axi_out_5_AR.valid" *)output m_axi_out_5_ARVALID;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [63:0] m_axi_out_5_AWADDR;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [1:0] m_axi_out_5_AWBURST;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [3:0] m_axi_out_5_AWCACHE;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [0:0] m_axi_out_5_AWID;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [7:0] m_axi_out_5_AWLEN;
  (* RS_HS = "m_axi_out_5_AW.data" *)output m_axi_out_5_AWLOCK;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [2:0] m_axi_out_5_AWPROT;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [3:0] m_axi_out_5_AWQOS;
  (* RS_HS = "m_axi_out_5_AW.ready" *)input m_axi_out_5_AWREADY;
  (* RS_HS = "m_axi_out_5_AW.data" *)output [2:0] m_axi_out_5_AWSIZE;
  (* RS_HS = "m_axi_out_5_AW.valid" *)output m_axi_out_5_AWVALID;
  (* RS_HS = "m_axi_out_5_B.data" *)input [0:0] m_axi_out_5_BID;
  (* RS_HS = "m_axi_out_5_B.ready" *)output m_axi_out_5_BREADY;
  (* RS_HS = "m_axi_out_5_B.data" *)input [1:0] m_axi_out_5_BRESP;
  (* RS_HS = "m_axi_out_5_B.valid" *)input m_axi_out_5_BVALID;
  (* RS_HS = "m_axi_out_5_R.data" *)input [511:0] m_axi_out_5_RDATA;
  (* RS_HS = "m_axi_out_5_R.data" *)input [0:0] m_axi_out_5_RID;
  (* RS_HS = "m_axi_out_5_R.data" *)input m_axi_out_5_RLAST;
  (* RS_HS = "m_axi_out_5_R.ready" *)output m_axi_out_5_RREADY;
  (* RS_HS = "m_axi_out_5_R.data" *)input [1:0] m_axi_out_5_RRESP;
  (* RS_HS = "m_axi_out_5_R.valid" *)input m_axi_out_5_RVALID;
  (* RS_HS = "m_axi_out_5_W.data" *)output [511:0] m_axi_out_5_WDATA;
  (* RS_HS = "m_axi_out_5_W.data" *)output m_axi_out_5_WLAST;
  (* RS_HS = "m_axi_out_5_W.ready" *)input m_axi_out_5_WREADY;
  (* RS_HS = "m_axi_out_5_W.data" *)output [63:0] m_axi_out_5_WSTRB;
  (* RS_HS = "m_axi_out_5_W.valid" *)output m_axi_out_5_WVALID;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [63:0] m_axi_in_6_ARADDR;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [1:0] m_axi_in_6_ARBURST;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [3:0] m_axi_in_6_ARCACHE;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [0:0] m_axi_in_6_ARID;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [7:0] m_axi_in_6_ARLEN;
  (* RS_HS = "m_axi_in_6_AR.data" *)output m_axi_in_6_ARLOCK;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [2:0] m_axi_in_6_ARPROT;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [3:0] m_axi_in_6_ARQOS;
  (* RS_HS = "m_axi_in_6_AR.ready" *)input m_axi_in_6_ARREADY;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [2:0] m_axi_in_6_ARSIZE;
  (* RS_HS = "m_axi_in_6_AR.valid" *)output m_axi_in_6_ARVALID;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [63:0] m_axi_in_6_AWADDR;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [1:0] m_axi_in_6_AWBURST;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [3:0] m_axi_in_6_AWCACHE;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [0:0] m_axi_in_6_AWID;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [7:0] m_axi_in_6_AWLEN;
  (* RS_HS = "m_axi_in_6_AW.data" *)output m_axi_in_6_AWLOCK;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [2:0] m_axi_in_6_AWPROT;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [3:0] m_axi_in_6_AWQOS;
  (* RS_HS = "m_axi_in_6_AW.ready" *)input m_axi_in_6_AWREADY;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [2:0] m_axi_in_6_AWSIZE;
  (* RS_HS = "m_axi_in_6_AW.valid" *)output m_axi_in_6_AWVALID;
  (* RS_HS = "m_axi_in_6_B.data" *)input [0:0] m_axi_in_6_BID;
  (* RS_HS = "m_axi_in_6_B.ready" *)output m_axi_in_6_BREADY;
  (* RS_HS = "m_axi_in_6_B.data" *)input [1:0] m_axi_in_6_BRESP;
  (* RS_HS = "m_axi_in_6_B.valid" *)input m_axi_in_6_BVALID;
  (* RS_HS = "m_axi_in_6_R.data" *)input [511:0] m_axi_in_6_RDATA;
  (* RS_HS = "m_axi_in_6_R.data" *)input [0:0] m_axi_in_6_RID;
  (* RS_HS = "m_axi_in_6_R.data" *)input m_axi_in_6_RLAST;
  (* RS_HS = "m_axi_in_6_R.ready" *)output m_axi_in_6_RREADY;
  (* RS_HS = "m_axi_in_6_R.data" *)input [1:0] m_axi_in_6_RRESP;
  (* RS_HS = "m_axi_in_6_R.valid" *)input m_axi_in_6_RVALID;
  (* RS_HS = "m_axi_in_6_W.data" *)output [511:0] m_axi_in_6_WDATA;
  (* RS_HS = "m_axi_in_6_W.data" *)output m_axi_in_6_WLAST;
  (* RS_HS = "m_axi_in_6_W.ready" *)input m_axi_in_6_WREADY;
  (* RS_HS = "m_axi_in_6_W.data" *)output [63:0] m_axi_in_6_WSTRB;
  (* RS_HS = "m_axi_in_6_W.valid" *)output m_axi_in_6_WVALID;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [63:0] m_axi_out_6_ARADDR;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [1:0] m_axi_out_6_ARBURST;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [3:0] m_axi_out_6_ARCACHE;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [0:0] m_axi_out_6_ARID;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [7:0] m_axi_out_6_ARLEN;
  (* RS_HS = "m_axi_out_6_AR.data" *)output m_axi_out_6_ARLOCK;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [2:0] m_axi_out_6_ARPROT;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [3:0] m_axi_out_6_ARQOS;
  (* RS_HS = "m_axi_out_6_AR.ready" *)input m_axi_out_6_ARREADY;
  (* RS_HS = "m_axi_out_6_AR.data" *)output [2:0] m_axi_out_6_ARSIZE;
  (* RS_HS = "m_axi_out_6_AR.valid" *)output m_axi_out_6_ARVALID;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [63:0] m_axi_out_6_AWADDR;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [1:0] m_axi_out_6_AWBURST;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [3:0] m_axi_out_6_AWCACHE;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [0:0] m_axi_out_6_AWID;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [7:0] m_axi_out_6_AWLEN;
  (* RS_HS = "m_axi_out_6_AW.data" *)output m_axi_out_6_AWLOCK;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [2:0] m_axi_out_6_AWPROT;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [3:0] m_axi_out_6_AWQOS;
  (* RS_HS = "m_axi_out_6_AW.ready" *)input m_axi_out_6_AWREADY;
  (* RS_HS = "m_axi_out_6_AW.data" *)output [2:0] m_axi_out_6_AWSIZE;
  (* RS_HS = "m_axi_out_6_AW.valid" *)output m_axi_out_6_AWVALID;
  (* RS_HS = "m_axi_out_6_B.data" *)input [0:0] m_axi_out_6_BID;
  (* RS_HS = "m_axi_out_6_B.ready" *)output m_axi_out_6_BREADY;
  (* RS_HS = "m_axi_out_6_B.data" *)input [1:0] m_axi_out_6_BRESP;
  (* RS_HS = "m_axi_out_6_B.valid" *)input m_axi_out_6_BVALID;
  (* RS_HS = "m_axi_out_6_R.data" *)input [511:0] m_axi_out_6_RDATA;
  (* RS_HS = "m_axi_out_6_R.data" *)input [0:0] m_axi_out_6_RID;
  (* RS_HS = "m_axi_out_6_R.data" *)input m_axi_out_6_RLAST;
  (* RS_HS = "m_axi_out_6_R.ready" *)output m_axi_out_6_RREADY;
  (* RS_HS = "m_axi_out_6_R.data" *)input [1:0] m_axi_out_6_RRESP;
  (* RS_HS = "m_axi_out_6_R.valid" *)input m_axi_out_6_RVALID;
  (* RS_HS = "m_axi_out_6_W.data" *)output [511:0] m_axi_out_6_WDATA;
  (* RS_HS = "m_axi_out_6_W.data" *)output m_axi_out_6_WLAST;
  (* RS_HS = "m_axi_out_6_W.ready" *)input m_axi_out_6_WREADY;
  (* RS_HS = "m_axi_out_6_W.data" *)output [63:0] m_axi_out_6_WSTRB;
  (* RS_HS = "m_axi_out_6_W.valid" *)output m_axi_out_6_WVALID;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [63:0] m_axi_in_7_ARADDR;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [1:0] m_axi_in_7_ARBURST;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [3:0] m_axi_in_7_ARCACHE;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [0:0] m_axi_in_7_ARID;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [7:0] m_axi_in_7_ARLEN;
  (* RS_HS = "m_axi_in_7_AR.data" *)output m_axi_in_7_ARLOCK;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [2:0] m_axi_in_7_ARPROT;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [3:0] m_axi_in_7_ARQOS;
  (* RS_HS = "m_axi_in_7_AR.ready" *)input m_axi_in_7_ARREADY;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [2:0] m_axi_in_7_ARSIZE;
  (* RS_HS = "m_axi_in_7_AR.valid" *)output m_axi_in_7_ARVALID;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [63:0] m_axi_in_7_AWADDR;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [1:0] m_axi_in_7_AWBURST;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [3:0] m_axi_in_7_AWCACHE;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [0:0] m_axi_in_7_AWID;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [7:0] m_axi_in_7_AWLEN;
  (* RS_HS = "m_axi_in_7_AW.data" *)output m_axi_in_7_AWLOCK;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [2:0] m_axi_in_7_AWPROT;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [3:0] m_axi_in_7_AWQOS;
  (* RS_HS = "m_axi_in_7_AW.ready" *)input m_axi_in_7_AWREADY;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [2:0] m_axi_in_7_AWSIZE;
  (* RS_HS = "m_axi_in_7_AW.valid" *)output m_axi_in_7_AWVALID;
  (* RS_HS = "m_axi_in_7_B.data" *)input [0:0] m_axi_in_7_BID;
  (* RS_HS = "m_axi_in_7_B.ready" *)output m_axi_in_7_BREADY;
  (* RS_HS = "m_axi_in_7_B.data" *)input [1:0] m_axi_in_7_BRESP;
  (* RS_HS = "m_axi_in_7_B.valid" *)input m_axi_in_7_BVALID;
  (* RS_HS = "m_axi_in_7_R.data" *)input [511:0] m_axi_in_7_RDATA;
  (* RS_HS = "m_axi_in_7_R.data" *)input [0:0] m_axi_in_7_RID;
  (* RS_HS = "m_axi_in_7_R.data" *)input m_axi_in_7_RLAST;
  (* RS_HS = "m_axi_in_7_R.ready" *)output m_axi_in_7_RREADY;
  (* RS_HS = "m_axi_in_7_R.data" *)input [1:0] m_axi_in_7_RRESP;
  (* RS_HS = "m_axi_in_7_R.valid" *)input m_axi_in_7_RVALID;
  (* RS_HS = "m_axi_in_7_W.data" *)output [511:0] m_axi_in_7_WDATA;
  (* RS_HS = "m_axi_in_7_W.data" *)output m_axi_in_7_WLAST;
  (* RS_HS = "m_axi_in_7_W.ready" *)input m_axi_in_7_WREADY;
  (* RS_HS = "m_axi_in_7_W.data" *)output [63:0] m_axi_in_7_WSTRB;
  (* RS_HS = "m_axi_in_7_W.valid" *)output m_axi_in_7_WVALID;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [63:0] m_axi_out_7_ARADDR;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [1:0] m_axi_out_7_ARBURST;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [3:0] m_axi_out_7_ARCACHE;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [0:0] m_axi_out_7_ARID;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [7:0] m_axi_out_7_ARLEN;
  (* RS_HS = "m_axi_out_7_AR.data" *)output m_axi_out_7_ARLOCK;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [2:0] m_axi_out_7_ARPROT;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [3:0] m_axi_out_7_ARQOS;
  (* RS_HS = "m_axi_out_7_AR.ready" *)input m_axi_out_7_ARREADY;
  (* RS_HS = "m_axi_out_7_AR.data" *)output [2:0] m_axi_out_7_ARSIZE;
  (* RS_HS = "m_axi_out_7_AR.valid" *)output m_axi_out_7_ARVALID;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [63:0] m_axi_out_7_AWADDR;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [1:0] m_axi_out_7_AWBURST;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [3:0] m_axi_out_7_AWCACHE;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [0:0] m_axi_out_7_AWID;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [7:0] m_axi_out_7_AWLEN;
  (* RS_HS = "m_axi_out_7_AW.data" *)output m_axi_out_7_AWLOCK;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [2:0] m_axi_out_7_AWPROT;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [3:0] m_axi_out_7_AWQOS;
  (* RS_HS = "m_axi_out_7_AW.ready" *)input m_axi_out_7_AWREADY;
  (* RS_HS = "m_axi_out_7_AW.data" *)output [2:0] m_axi_out_7_AWSIZE;
  (* RS_HS = "m_axi_out_7_AW.valid" *)output m_axi_out_7_AWVALID;
  (* RS_HS = "m_axi_out_7_B.data" *)input [0:0] m_axi_out_7_BID;
  (* RS_HS = "m_axi_out_7_B.ready" *)output m_axi_out_7_BREADY;
  (* RS_HS = "m_axi_out_7_B.data" *)input [1:0] m_axi_out_7_BRESP;
  (* RS_HS = "m_axi_out_7_B.valid" *)input m_axi_out_7_BVALID;
  (* RS_HS = "m_axi_out_7_R.data" *)input [511:0] m_axi_out_7_RDATA;
  (* RS_HS = "m_axi_out_7_R.data" *)input [0:0] m_axi_out_7_RID;
  (* RS_HS = "m_axi_out_7_R.data" *)input m_axi_out_7_RLAST;
  (* RS_HS = "m_axi_out_7_R.ready" *)output m_axi_out_7_RREADY;
  (* RS_HS = "m_axi_out_7_R.data" *)input [1:0] m_axi_out_7_RRESP;
  (* RS_HS = "m_axi_out_7_R.valid" *)input m_axi_out_7_RVALID;
  (* RS_HS = "m_axi_out_7_W.data" *)output [511:0] m_axi_out_7_WDATA;
  (* RS_HS = "m_axi_out_7_W.data" *)output m_axi_out_7_WLAST;
  (* RS_HS = "m_axi_out_7_W.ready" *)input m_axi_out_7_WREADY;
  (* RS_HS = "m_axi_out_7_W.data" *)output [63:0] m_axi_out_7_WSTRB;
  (* RS_HS = "m_axi_out_7_W.valid" *)output m_axi_out_7_WVALID;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [63:0] m_axi_in_8_ARADDR;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [1:0] m_axi_in_8_ARBURST;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [3:0] m_axi_in_8_ARCACHE;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [0:0] m_axi_in_8_ARID;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [7:0] m_axi_in_8_ARLEN;
  (* RS_HS = "m_axi_in_8_AR.data" *)output m_axi_in_8_ARLOCK;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [2:0] m_axi_in_8_ARPROT;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [3:0] m_axi_in_8_ARQOS;
  (* RS_HS = "m_axi_in_8_AR.ready" *)input m_axi_in_8_ARREADY;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [2:0] m_axi_in_8_ARSIZE;
  (* RS_HS = "m_axi_in_8_AR.valid" *)output m_axi_in_8_ARVALID;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [63:0] m_axi_in_8_AWADDR;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [1:0] m_axi_in_8_AWBURST;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [3:0] m_axi_in_8_AWCACHE;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [0:0] m_axi_in_8_AWID;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [7:0] m_axi_in_8_AWLEN;
  (* RS_HS = "m_axi_in_8_AW.data" *)output m_axi_in_8_AWLOCK;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [2:0] m_axi_in_8_AWPROT;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [3:0] m_axi_in_8_AWQOS;
  (* RS_HS = "m_axi_in_8_AW.ready" *)input m_axi_in_8_AWREADY;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [2:0] m_axi_in_8_AWSIZE;
  (* RS_HS = "m_axi_in_8_AW.valid" *)output m_axi_in_8_AWVALID;
  (* RS_HS = "m_axi_in_8_B.data" *)input [0:0] m_axi_in_8_BID;
  (* RS_HS = "m_axi_in_8_B.ready" *)output m_axi_in_8_BREADY;
  (* RS_HS = "m_axi_in_8_B.data" *)input [1:0] m_axi_in_8_BRESP;
  (* RS_HS = "m_axi_in_8_B.valid" *)input m_axi_in_8_BVALID;
  (* RS_HS = "m_axi_in_8_R.data" *)input [511:0] m_axi_in_8_RDATA;
  (* RS_HS = "m_axi_in_8_R.data" *)input [0:0] m_axi_in_8_RID;
  (* RS_HS = "m_axi_in_8_R.data" *)input m_axi_in_8_RLAST;
  (* RS_HS = "m_axi_in_8_R.ready" *)output m_axi_in_8_RREADY;
  (* RS_HS = "m_axi_in_8_R.data" *)input [1:0] m_axi_in_8_RRESP;
  (* RS_HS = "m_axi_in_8_R.valid" *)input m_axi_in_8_RVALID;
  (* RS_HS = "m_axi_in_8_W.data" *)output [511:0] m_axi_in_8_WDATA;
  (* RS_HS = "m_axi_in_8_W.data" *)output m_axi_in_8_WLAST;
  (* RS_HS = "m_axi_in_8_W.ready" *)input m_axi_in_8_WREADY;
  (* RS_HS = "m_axi_in_8_W.data" *)output [63:0] m_axi_in_8_WSTRB;
  (* RS_HS = "m_axi_in_8_W.valid" *)output m_axi_in_8_WVALID;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [63:0] m_axi_out_8_ARADDR;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [1:0] m_axi_out_8_ARBURST;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [3:0] m_axi_out_8_ARCACHE;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [0:0] m_axi_out_8_ARID;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [7:0] m_axi_out_8_ARLEN;
  (* RS_HS = "m_axi_out_8_AR.data" *)output m_axi_out_8_ARLOCK;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [2:0] m_axi_out_8_ARPROT;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [3:0] m_axi_out_8_ARQOS;
  (* RS_HS = "m_axi_out_8_AR.ready" *)input m_axi_out_8_ARREADY;
  (* RS_HS = "m_axi_out_8_AR.data" *)output [2:0] m_axi_out_8_ARSIZE;
  (* RS_HS = "m_axi_out_8_AR.valid" *)output m_axi_out_8_ARVALID;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [63:0] m_axi_out_8_AWADDR;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [1:0] m_axi_out_8_AWBURST;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [3:0] m_axi_out_8_AWCACHE;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [0:0] m_axi_out_8_AWID;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [7:0] m_axi_out_8_AWLEN;
  (* RS_HS = "m_axi_out_8_AW.data" *)output m_axi_out_8_AWLOCK;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [2:0] m_axi_out_8_AWPROT;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [3:0] m_axi_out_8_AWQOS;
  (* RS_HS = "m_axi_out_8_AW.ready" *)input m_axi_out_8_AWREADY;
  (* RS_HS = "m_axi_out_8_AW.data" *)output [2:0] m_axi_out_8_AWSIZE;
  (* RS_HS = "m_axi_out_8_AW.valid" *)output m_axi_out_8_AWVALID;
  (* RS_HS = "m_axi_out_8_B.data" *)input [0:0] m_axi_out_8_BID;
  (* RS_HS = "m_axi_out_8_B.ready" *)output m_axi_out_8_BREADY;
  (* RS_HS = "m_axi_out_8_B.data" *)input [1:0] m_axi_out_8_BRESP;
  (* RS_HS = "m_axi_out_8_B.valid" *)input m_axi_out_8_BVALID;
  (* RS_HS = "m_axi_out_8_R.data" *)input [511:0] m_axi_out_8_RDATA;
  (* RS_HS = "m_axi_out_8_R.data" *)input [0:0] m_axi_out_8_RID;
  (* RS_HS = "m_axi_out_8_R.data" *)input m_axi_out_8_RLAST;
  (* RS_HS = "m_axi_out_8_R.ready" *)output m_axi_out_8_RREADY;
  (* RS_HS = "m_axi_out_8_R.data" *)input [1:0] m_axi_out_8_RRESP;
  (* RS_HS = "m_axi_out_8_R.valid" *)input m_axi_out_8_RVALID;
  (* RS_HS = "m_axi_out_8_W.data" *)output [511:0] m_axi_out_8_WDATA;
  (* RS_HS = "m_axi_out_8_W.data" *)output m_axi_out_8_WLAST;
  (* RS_HS = "m_axi_out_8_W.ready" *)input m_axi_out_8_WREADY;
  (* RS_HS = "m_axi_out_8_W.data" *)output [63:0] m_axi_out_8_WSTRB;
  (* RS_HS = "m_axi_out_8_W.valid" *)output m_axi_out_8_WVALID;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [63:0] m_axi_in_9_ARADDR;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [1:0] m_axi_in_9_ARBURST;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [3:0] m_axi_in_9_ARCACHE;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [0:0] m_axi_in_9_ARID;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [7:0] m_axi_in_9_ARLEN;
  (* RS_HS = "m_axi_in_9_AR.data" *)output m_axi_in_9_ARLOCK;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [2:0] m_axi_in_9_ARPROT;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [3:0] m_axi_in_9_ARQOS;
  (* RS_HS = "m_axi_in_9_AR.ready" *)input m_axi_in_9_ARREADY;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [2:0] m_axi_in_9_ARSIZE;
  (* RS_HS = "m_axi_in_9_AR.valid" *)output m_axi_in_9_ARVALID;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [63:0] m_axi_in_9_AWADDR;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [1:0] m_axi_in_9_AWBURST;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [3:0] m_axi_in_9_AWCACHE;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [0:0] m_axi_in_9_AWID;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [7:0] m_axi_in_9_AWLEN;
  (* RS_HS = "m_axi_in_9_AW.data" *)output m_axi_in_9_AWLOCK;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [2:0] m_axi_in_9_AWPROT;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [3:0] m_axi_in_9_AWQOS;
  (* RS_HS = "m_axi_in_9_AW.ready" *)input m_axi_in_9_AWREADY;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [2:0] m_axi_in_9_AWSIZE;
  (* RS_HS = "m_axi_in_9_AW.valid" *)output m_axi_in_9_AWVALID;
  (* RS_HS = "m_axi_in_9_B.data" *)input [0:0] m_axi_in_9_BID;
  (* RS_HS = "m_axi_in_9_B.ready" *)output m_axi_in_9_BREADY;
  (* RS_HS = "m_axi_in_9_B.data" *)input [1:0] m_axi_in_9_BRESP;
  (* RS_HS = "m_axi_in_9_B.valid" *)input m_axi_in_9_BVALID;
  (* RS_HS = "m_axi_in_9_R.data" *)input [511:0] m_axi_in_9_RDATA;
  (* RS_HS = "m_axi_in_9_R.data" *)input [0:0] m_axi_in_9_RID;
  (* RS_HS = "m_axi_in_9_R.data" *)input m_axi_in_9_RLAST;
  (* RS_HS = "m_axi_in_9_R.ready" *)output m_axi_in_9_RREADY;
  (* RS_HS = "m_axi_in_9_R.data" *)input [1:0] m_axi_in_9_RRESP;
  (* RS_HS = "m_axi_in_9_R.valid" *)input m_axi_in_9_RVALID;
  (* RS_HS = "m_axi_in_9_W.data" *)output [511:0] m_axi_in_9_WDATA;
  (* RS_HS = "m_axi_in_9_W.data" *)output m_axi_in_9_WLAST;
  (* RS_HS = "m_axi_in_9_W.ready" *)input m_axi_in_9_WREADY;
  (* RS_HS = "m_axi_in_9_W.data" *)output [63:0] m_axi_in_9_WSTRB;
  (* RS_HS = "m_axi_in_9_W.valid" *)output m_axi_in_9_WVALID;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [63:0] m_axi_out_9_ARADDR;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [1:0] m_axi_out_9_ARBURST;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [3:0] m_axi_out_9_ARCACHE;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [0:0] m_axi_out_9_ARID;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [7:0] m_axi_out_9_ARLEN;
  (* RS_HS = "m_axi_out_9_AR.data" *)output m_axi_out_9_ARLOCK;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [2:0] m_axi_out_9_ARPROT;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [3:0] m_axi_out_9_ARQOS;
  (* RS_HS = "m_axi_out_9_AR.ready" *)input m_axi_out_9_ARREADY;
  (* RS_HS = "m_axi_out_9_AR.data" *)output [2:0] m_axi_out_9_ARSIZE;
  (* RS_HS = "m_axi_out_9_AR.valid" *)output m_axi_out_9_ARVALID;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [63:0] m_axi_out_9_AWADDR;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [1:0] m_axi_out_9_AWBURST;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [3:0] m_axi_out_9_AWCACHE;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [0:0] m_axi_out_9_AWID;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [7:0] m_axi_out_9_AWLEN;
  (* RS_HS = "m_axi_out_9_AW.data" *)output m_axi_out_9_AWLOCK;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [2:0] m_axi_out_9_AWPROT;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [3:0] m_axi_out_9_AWQOS;
  (* RS_HS = "m_axi_out_9_AW.ready" *)input m_axi_out_9_AWREADY;
  (* RS_HS = "m_axi_out_9_AW.data" *)output [2:0] m_axi_out_9_AWSIZE;
  (* RS_HS = "m_axi_out_9_AW.valid" *)output m_axi_out_9_AWVALID;
  (* RS_HS = "m_axi_out_9_B.data" *)input [0:0] m_axi_out_9_BID;
  (* RS_HS = "m_axi_out_9_B.ready" *)output m_axi_out_9_BREADY;
  (* RS_HS = "m_axi_out_9_B.data" *)input [1:0] m_axi_out_9_BRESP;
  (* RS_HS = "m_axi_out_9_B.valid" *)input m_axi_out_9_BVALID;
  (* RS_HS = "m_axi_out_9_R.data" *)input [511:0] m_axi_out_9_RDATA;
  (* RS_HS = "m_axi_out_9_R.data" *)input [0:0] m_axi_out_9_RID;
  (* RS_HS = "m_axi_out_9_R.data" *)input m_axi_out_9_RLAST;
  (* RS_HS = "m_axi_out_9_R.ready" *)output m_axi_out_9_RREADY;
  (* RS_HS = "m_axi_out_9_R.data" *)input [1:0] m_axi_out_9_RRESP;
  (* RS_HS = "m_axi_out_9_R.valid" *)input m_axi_out_9_RVALID;
  (* RS_HS = "m_axi_out_9_W.data" *)output [511:0] m_axi_out_9_WDATA;
  (* RS_HS = "m_axi_out_9_W.data" *)output m_axi_out_9_WLAST;
  (* RS_HS = "m_axi_out_9_W.ready" *)input m_axi_out_9_WREADY;
  (* RS_HS = "m_axi_out_9_W.data" *)output [63:0] m_axi_out_9_WSTRB;
  (* RS_HS = "m_axi_out_9_W.valid" *)output m_axi_out_9_WVALID;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [63:0] m_axi_in_10_ARADDR;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [1:0] m_axi_in_10_ARBURST;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [3:0] m_axi_in_10_ARCACHE;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [0:0] m_axi_in_10_ARID;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [7:0] m_axi_in_10_ARLEN;
  (* RS_HS = "m_axi_in_10_AR.data" *)output m_axi_in_10_ARLOCK;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [2:0] m_axi_in_10_ARPROT;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [3:0] m_axi_in_10_ARQOS;
  (* RS_HS = "m_axi_in_10_AR.ready" *)input m_axi_in_10_ARREADY;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [2:0] m_axi_in_10_ARSIZE;
  (* RS_HS = "m_axi_in_10_AR.valid" *)output m_axi_in_10_ARVALID;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [63:0] m_axi_in_10_AWADDR;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [1:0] m_axi_in_10_AWBURST;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [3:0] m_axi_in_10_AWCACHE;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [0:0] m_axi_in_10_AWID;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [7:0] m_axi_in_10_AWLEN;
  (* RS_HS = "m_axi_in_10_AW.data" *)output m_axi_in_10_AWLOCK;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [2:0] m_axi_in_10_AWPROT;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [3:0] m_axi_in_10_AWQOS;
  (* RS_HS = "m_axi_in_10_AW.ready" *)input m_axi_in_10_AWREADY;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [2:0] m_axi_in_10_AWSIZE;
  (* RS_HS = "m_axi_in_10_AW.valid" *)output m_axi_in_10_AWVALID;
  (* RS_HS = "m_axi_in_10_B.data" *)input [0:0] m_axi_in_10_BID;
  (* RS_HS = "m_axi_in_10_B.ready" *)output m_axi_in_10_BREADY;
  (* RS_HS = "m_axi_in_10_B.data" *)input [1:0] m_axi_in_10_BRESP;
  (* RS_HS = "m_axi_in_10_B.valid" *)input m_axi_in_10_BVALID;
  (* RS_HS = "m_axi_in_10_R.data" *)input [511:0] m_axi_in_10_RDATA;
  (* RS_HS = "m_axi_in_10_R.data" *)input [0:0] m_axi_in_10_RID;
  (* RS_HS = "m_axi_in_10_R.data" *)input m_axi_in_10_RLAST;
  (* RS_HS = "m_axi_in_10_R.ready" *)output m_axi_in_10_RREADY;
  (* RS_HS = "m_axi_in_10_R.data" *)input [1:0] m_axi_in_10_RRESP;
  (* RS_HS = "m_axi_in_10_R.valid" *)input m_axi_in_10_RVALID;
  (* RS_HS = "m_axi_in_10_W.data" *)output [511:0] m_axi_in_10_WDATA;
  (* RS_HS = "m_axi_in_10_W.data" *)output m_axi_in_10_WLAST;
  (* RS_HS = "m_axi_in_10_W.ready" *)input m_axi_in_10_WREADY;
  (* RS_HS = "m_axi_in_10_W.data" *)output [63:0] m_axi_in_10_WSTRB;
  (* RS_HS = "m_axi_in_10_W.valid" *)output m_axi_in_10_WVALID;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [63:0] m_axi_out_10_ARADDR;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [1:0] m_axi_out_10_ARBURST;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [3:0] m_axi_out_10_ARCACHE;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [0:0] m_axi_out_10_ARID;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [7:0] m_axi_out_10_ARLEN;
  (* RS_HS = "m_axi_out_10_AR.data" *)output m_axi_out_10_ARLOCK;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [2:0] m_axi_out_10_ARPROT;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [3:0] m_axi_out_10_ARQOS;
  (* RS_HS = "m_axi_out_10_AR.ready" *)input m_axi_out_10_ARREADY;
  (* RS_HS = "m_axi_out_10_AR.data" *)output [2:0] m_axi_out_10_ARSIZE;
  (* RS_HS = "m_axi_out_10_AR.valid" *)output m_axi_out_10_ARVALID;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [63:0] m_axi_out_10_AWADDR;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [1:0] m_axi_out_10_AWBURST;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [3:0] m_axi_out_10_AWCACHE;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [0:0] m_axi_out_10_AWID;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [7:0] m_axi_out_10_AWLEN;
  (* RS_HS = "m_axi_out_10_AW.data" *)output m_axi_out_10_AWLOCK;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [2:0] m_axi_out_10_AWPROT;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [3:0] m_axi_out_10_AWQOS;
  (* RS_HS = "m_axi_out_10_AW.ready" *)input m_axi_out_10_AWREADY;
  (* RS_HS = "m_axi_out_10_AW.data" *)output [2:0] m_axi_out_10_AWSIZE;
  (* RS_HS = "m_axi_out_10_AW.valid" *)output m_axi_out_10_AWVALID;
  (* RS_HS = "m_axi_out_10_B.data" *)input [0:0] m_axi_out_10_BID;
  (* RS_HS = "m_axi_out_10_B.ready" *)output m_axi_out_10_BREADY;
  (* RS_HS = "m_axi_out_10_B.data" *)input [1:0] m_axi_out_10_BRESP;
  (* RS_HS = "m_axi_out_10_B.valid" *)input m_axi_out_10_BVALID;
  (* RS_HS = "m_axi_out_10_R.data" *)input [511:0] m_axi_out_10_RDATA;
  (* RS_HS = "m_axi_out_10_R.data" *)input [0:0] m_axi_out_10_RID;
  (* RS_HS = "m_axi_out_10_R.data" *)input m_axi_out_10_RLAST;
  (* RS_HS = "m_axi_out_10_R.ready" *)output m_axi_out_10_RREADY;
  (* RS_HS = "m_axi_out_10_R.data" *)input [1:0] m_axi_out_10_RRESP;
  (* RS_HS = "m_axi_out_10_R.valid" *)input m_axi_out_10_RVALID;
  (* RS_HS = "m_axi_out_10_W.data" *)output [511:0] m_axi_out_10_WDATA;
  (* RS_HS = "m_axi_out_10_W.data" *)output m_axi_out_10_WLAST;
  (* RS_HS = "m_axi_out_10_W.ready" *)input m_axi_out_10_WREADY;
  (* RS_HS = "m_axi_out_10_W.data" *)output [63:0] m_axi_out_10_WSTRB;
  (* RS_HS = "m_axi_out_10_W.valid" *)output m_axi_out_10_WVALID;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [63:0] m_axi_in_11_ARADDR;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [1:0] m_axi_in_11_ARBURST;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [3:0] m_axi_in_11_ARCACHE;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [0:0] m_axi_in_11_ARID;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [7:0] m_axi_in_11_ARLEN;
  (* RS_HS = "m_axi_in_11_AR.data" *)output m_axi_in_11_ARLOCK;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [2:0] m_axi_in_11_ARPROT;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [3:0] m_axi_in_11_ARQOS;
  (* RS_HS = "m_axi_in_11_AR.ready" *)input m_axi_in_11_ARREADY;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [2:0] m_axi_in_11_ARSIZE;
  (* RS_HS = "m_axi_in_11_AR.valid" *)output m_axi_in_11_ARVALID;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [63:0] m_axi_in_11_AWADDR;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [1:0] m_axi_in_11_AWBURST;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [3:0] m_axi_in_11_AWCACHE;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [0:0] m_axi_in_11_AWID;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [7:0] m_axi_in_11_AWLEN;
  (* RS_HS = "m_axi_in_11_AW.data" *)output m_axi_in_11_AWLOCK;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [2:0] m_axi_in_11_AWPROT;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [3:0] m_axi_in_11_AWQOS;
  (* RS_HS = "m_axi_in_11_AW.ready" *)input m_axi_in_11_AWREADY;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [2:0] m_axi_in_11_AWSIZE;
  (* RS_HS = "m_axi_in_11_AW.valid" *)output m_axi_in_11_AWVALID;
  (* RS_HS = "m_axi_in_11_B.data" *)input [0:0] m_axi_in_11_BID;
  (* RS_HS = "m_axi_in_11_B.ready" *)output m_axi_in_11_BREADY;
  (* RS_HS = "m_axi_in_11_B.data" *)input [1:0] m_axi_in_11_BRESP;
  (* RS_HS = "m_axi_in_11_B.valid" *)input m_axi_in_11_BVALID;
  (* RS_HS = "m_axi_in_11_R.data" *)input [511:0] m_axi_in_11_RDATA;
  (* RS_HS = "m_axi_in_11_R.data" *)input [0:0] m_axi_in_11_RID;
  (* RS_HS = "m_axi_in_11_R.data" *)input m_axi_in_11_RLAST;
  (* RS_HS = "m_axi_in_11_R.ready" *)output m_axi_in_11_RREADY;
  (* RS_HS = "m_axi_in_11_R.data" *)input [1:0] m_axi_in_11_RRESP;
  (* RS_HS = "m_axi_in_11_R.valid" *)input m_axi_in_11_RVALID;
  (* RS_HS = "m_axi_in_11_W.data" *)output [511:0] m_axi_in_11_WDATA;
  (* RS_HS = "m_axi_in_11_W.data" *)output m_axi_in_11_WLAST;
  (* RS_HS = "m_axi_in_11_W.ready" *)input m_axi_in_11_WREADY;
  (* RS_HS = "m_axi_in_11_W.data" *)output [63:0] m_axi_in_11_WSTRB;
  (* RS_HS = "m_axi_in_11_W.valid" *)output m_axi_in_11_WVALID;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [63:0] m_axi_out_11_ARADDR;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [1:0] m_axi_out_11_ARBURST;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [3:0] m_axi_out_11_ARCACHE;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [0:0] m_axi_out_11_ARID;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [7:0] m_axi_out_11_ARLEN;
  (* RS_HS = "m_axi_out_11_AR.data" *)output m_axi_out_11_ARLOCK;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [2:0] m_axi_out_11_ARPROT;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [3:0] m_axi_out_11_ARQOS;
  (* RS_HS = "m_axi_out_11_AR.ready" *)input m_axi_out_11_ARREADY;
  (* RS_HS = "m_axi_out_11_AR.data" *)output [2:0] m_axi_out_11_ARSIZE;
  (* RS_HS = "m_axi_out_11_AR.valid" *)output m_axi_out_11_ARVALID;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [63:0] m_axi_out_11_AWADDR;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [1:0] m_axi_out_11_AWBURST;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [3:0] m_axi_out_11_AWCACHE;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [0:0] m_axi_out_11_AWID;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [7:0] m_axi_out_11_AWLEN;
  (* RS_HS = "m_axi_out_11_AW.data" *)output m_axi_out_11_AWLOCK;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [2:0] m_axi_out_11_AWPROT;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [3:0] m_axi_out_11_AWQOS;
  (* RS_HS = "m_axi_out_11_AW.ready" *)input m_axi_out_11_AWREADY;
  (* RS_HS = "m_axi_out_11_AW.data" *)output [2:0] m_axi_out_11_AWSIZE;
  (* RS_HS = "m_axi_out_11_AW.valid" *)output m_axi_out_11_AWVALID;
  (* RS_HS = "m_axi_out_11_B.data" *)input [0:0] m_axi_out_11_BID;
  (* RS_HS = "m_axi_out_11_B.ready" *)output m_axi_out_11_BREADY;
  (* RS_HS = "m_axi_out_11_B.data" *)input [1:0] m_axi_out_11_BRESP;
  (* RS_HS = "m_axi_out_11_B.valid" *)input m_axi_out_11_BVALID;
  (* RS_HS = "m_axi_out_11_R.data" *)input [511:0] m_axi_out_11_RDATA;
  (* RS_HS = "m_axi_out_11_R.data" *)input [0:0] m_axi_out_11_RID;
  (* RS_HS = "m_axi_out_11_R.data" *)input m_axi_out_11_RLAST;
  (* RS_HS = "m_axi_out_11_R.ready" *)output m_axi_out_11_RREADY;
  (* RS_HS = "m_axi_out_11_R.data" *)input [1:0] m_axi_out_11_RRESP;
  (* RS_HS = "m_axi_out_11_R.valid" *)input m_axi_out_11_RVALID;
  (* RS_HS = "m_axi_out_11_W.data" *)output [511:0] m_axi_out_11_WDATA;
  (* RS_HS = "m_axi_out_11_W.data" *)output m_axi_out_11_WLAST;
  (* RS_HS = "m_axi_out_11_W.ready" *)input m_axi_out_11_WREADY;
  (* RS_HS = "m_axi_out_11_W.data" *)output [63:0] m_axi_out_11_WSTRB;
  (* RS_HS = "m_axi_out_11_W.valid" *)output m_axi_out_11_WVALID;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [63:0] m_axi_in_12_ARADDR;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [1:0] m_axi_in_12_ARBURST;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [3:0] m_axi_in_12_ARCACHE;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [0:0] m_axi_in_12_ARID;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [7:0] m_axi_in_12_ARLEN;
  (* RS_HS = "m_axi_in_12_AR.data" *)output m_axi_in_12_ARLOCK;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [2:0] m_axi_in_12_ARPROT;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [3:0] m_axi_in_12_ARQOS;
  (* RS_HS = "m_axi_in_12_AR.ready" *)input m_axi_in_12_ARREADY;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [2:0] m_axi_in_12_ARSIZE;
  (* RS_HS = "m_axi_in_12_AR.valid" *)output m_axi_in_12_ARVALID;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [63:0] m_axi_in_12_AWADDR;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [1:0] m_axi_in_12_AWBURST;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [3:0] m_axi_in_12_AWCACHE;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [0:0] m_axi_in_12_AWID;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [7:0] m_axi_in_12_AWLEN;
  (* RS_HS = "m_axi_in_12_AW.data" *)output m_axi_in_12_AWLOCK;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [2:0] m_axi_in_12_AWPROT;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [3:0] m_axi_in_12_AWQOS;
  (* RS_HS = "m_axi_in_12_AW.ready" *)input m_axi_in_12_AWREADY;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [2:0] m_axi_in_12_AWSIZE;
  (* RS_HS = "m_axi_in_12_AW.valid" *)output m_axi_in_12_AWVALID;
  (* RS_HS = "m_axi_in_12_B.data" *)input [0:0] m_axi_in_12_BID;
  (* RS_HS = "m_axi_in_12_B.ready" *)output m_axi_in_12_BREADY;
  (* RS_HS = "m_axi_in_12_B.data" *)input [1:0] m_axi_in_12_BRESP;
  (* RS_HS = "m_axi_in_12_B.valid" *)input m_axi_in_12_BVALID;
  (* RS_HS = "m_axi_in_12_R.data" *)input [511:0] m_axi_in_12_RDATA;
  (* RS_HS = "m_axi_in_12_R.data" *)input [0:0] m_axi_in_12_RID;
  (* RS_HS = "m_axi_in_12_R.data" *)input m_axi_in_12_RLAST;
  (* RS_HS = "m_axi_in_12_R.ready" *)output m_axi_in_12_RREADY;
  (* RS_HS = "m_axi_in_12_R.data" *)input [1:0] m_axi_in_12_RRESP;
  (* RS_HS = "m_axi_in_12_R.valid" *)input m_axi_in_12_RVALID;
  (* RS_HS = "m_axi_in_12_W.data" *)output [511:0] m_axi_in_12_WDATA;
  (* RS_HS = "m_axi_in_12_W.data" *)output m_axi_in_12_WLAST;
  (* RS_HS = "m_axi_in_12_W.ready" *)input m_axi_in_12_WREADY;
  (* RS_HS = "m_axi_in_12_W.data" *)output [63:0] m_axi_in_12_WSTRB;
  (* RS_HS = "m_axi_in_12_W.valid" *)output m_axi_in_12_WVALID;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [63:0] m_axi_out_12_ARADDR;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [1:0] m_axi_out_12_ARBURST;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [3:0] m_axi_out_12_ARCACHE;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [0:0] m_axi_out_12_ARID;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [7:0] m_axi_out_12_ARLEN;
  (* RS_HS = "m_axi_out_12_AR.data" *)output m_axi_out_12_ARLOCK;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [2:0] m_axi_out_12_ARPROT;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [3:0] m_axi_out_12_ARQOS;
  (* RS_HS = "m_axi_out_12_AR.ready" *)input m_axi_out_12_ARREADY;
  (* RS_HS = "m_axi_out_12_AR.data" *)output [2:0] m_axi_out_12_ARSIZE;
  (* RS_HS = "m_axi_out_12_AR.valid" *)output m_axi_out_12_ARVALID;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [63:0] m_axi_out_12_AWADDR;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [1:0] m_axi_out_12_AWBURST;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [3:0] m_axi_out_12_AWCACHE;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [0:0] m_axi_out_12_AWID;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [7:0] m_axi_out_12_AWLEN;
  (* RS_HS = "m_axi_out_12_AW.data" *)output m_axi_out_12_AWLOCK;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [2:0] m_axi_out_12_AWPROT;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [3:0] m_axi_out_12_AWQOS;
  (* RS_HS = "m_axi_out_12_AW.ready" *)input m_axi_out_12_AWREADY;
  (* RS_HS = "m_axi_out_12_AW.data" *)output [2:0] m_axi_out_12_AWSIZE;
  (* RS_HS = "m_axi_out_12_AW.valid" *)output m_axi_out_12_AWVALID;
  (* RS_HS = "m_axi_out_12_B.data" *)input [0:0] m_axi_out_12_BID;
  (* RS_HS = "m_axi_out_12_B.ready" *)output m_axi_out_12_BREADY;
  (* RS_HS = "m_axi_out_12_B.data" *)input [1:0] m_axi_out_12_BRESP;
  (* RS_HS = "m_axi_out_12_B.valid" *)input m_axi_out_12_BVALID;
  (* RS_HS = "m_axi_out_12_R.data" *)input [511:0] m_axi_out_12_RDATA;
  (* RS_HS = "m_axi_out_12_R.data" *)input [0:0] m_axi_out_12_RID;
  (* RS_HS = "m_axi_out_12_R.data" *)input m_axi_out_12_RLAST;
  (* RS_HS = "m_axi_out_12_R.ready" *)output m_axi_out_12_RREADY;
  (* RS_HS = "m_axi_out_12_R.data" *)input [1:0] m_axi_out_12_RRESP;
  (* RS_HS = "m_axi_out_12_R.valid" *)input m_axi_out_12_RVALID;
  (* RS_HS = "m_axi_out_12_W.data" *)output [511:0] m_axi_out_12_WDATA;
  (* RS_HS = "m_axi_out_12_W.data" *)output m_axi_out_12_WLAST;
  (* RS_HS = "m_axi_out_12_W.ready" *)input m_axi_out_12_WREADY;
  (* RS_HS = "m_axi_out_12_W.data" *)output [63:0] m_axi_out_12_WSTRB;
  (* RS_HS = "m_axi_out_12_W.valid" *)output m_axi_out_12_WVALID;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [63:0] m_axi_in_13_ARADDR;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [1:0] m_axi_in_13_ARBURST;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [3:0] m_axi_in_13_ARCACHE;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [0:0] m_axi_in_13_ARID;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [7:0] m_axi_in_13_ARLEN;
  (* RS_HS = "m_axi_in_13_AR.data" *)output m_axi_in_13_ARLOCK;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [2:0] m_axi_in_13_ARPROT;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [3:0] m_axi_in_13_ARQOS;
  (* RS_HS = "m_axi_in_13_AR.ready" *)input m_axi_in_13_ARREADY;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [2:0] m_axi_in_13_ARSIZE;
  (* RS_HS = "m_axi_in_13_AR.valid" *)output m_axi_in_13_ARVALID;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [63:0] m_axi_in_13_AWADDR;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [1:0] m_axi_in_13_AWBURST;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [3:0] m_axi_in_13_AWCACHE;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [0:0] m_axi_in_13_AWID;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [7:0] m_axi_in_13_AWLEN;
  (* RS_HS = "m_axi_in_13_AW.data" *)output m_axi_in_13_AWLOCK;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [2:0] m_axi_in_13_AWPROT;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [3:0] m_axi_in_13_AWQOS;
  (* RS_HS = "m_axi_in_13_AW.ready" *)input m_axi_in_13_AWREADY;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [2:0] m_axi_in_13_AWSIZE;
  (* RS_HS = "m_axi_in_13_AW.valid" *)output m_axi_in_13_AWVALID;
  (* RS_HS = "m_axi_in_13_B.data" *)input [0:0] m_axi_in_13_BID;
  (* RS_HS = "m_axi_in_13_B.ready" *)output m_axi_in_13_BREADY;
  (* RS_HS = "m_axi_in_13_B.data" *)input [1:0] m_axi_in_13_BRESP;
  (* RS_HS = "m_axi_in_13_B.valid" *)input m_axi_in_13_BVALID;
  (* RS_HS = "m_axi_in_13_R.data" *)input [511:0] m_axi_in_13_RDATA;
  (* RS_HS = "m_axi_in_13_R.data" *)input [0:0] m_axi_in_13_RID;
  (* RS_HS = "m_axi_in_13_R.data" *)input m_axi_in_13_RLAST;
  (* RS_HS = "m_axi_in_13_R.ready" *)output m_axi_in_13_RREADY;
  (* RS_HS = "m_axi_in_13_R.data" *)input [1:0] m_axi_in_13_RRESP;
  (* RS_HS = "m_axi_in_13_R.valid" *)input m_axi_in_13_RVALID;
  (* RS_HS = "m_axi_in_13_W.data" *)output [511:0] m_axi_in_13_WDATA;
  (* RS_HS = "m_axi_in_13_W.data" *)output m_axi_in_13_WLAST;
  (* RS_HS = "m_axi_in_13_W.ready" *)input m_axi_in_13_WREADY;
  (* RS_HS = "m_axi_in_13_W.data" *)output [63:0] m_axi_in_13_WSTRB;
  (* RS_HS = "m_axi_in_13_W.valid" *)output m_axi_in_13_WVALID;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [63:0] m_axi_out_13_ARADDR;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [1:0] m_axi_out_13_ARBURST;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [3:0] m_axi_out_13_ARCACHE;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [0:0] m_axi_out_13_ARID;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [7:0] m_axi_out_13_ARLEN;
  (* RS_HS = "m_axi_out_13_AR.data" *)output m_axi_out_13_ARLOCK;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [2:0] m_axi_out_13_ARPROT;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [3:0] m_axi_out_13_ARQOS;
  (* RS_HS = "m_axi_out_13_AR.ready" *)input m_axi_out_13_ARREADY;
  (* RS_HS = "m_axi_out_13_AR.data" *)output [2:0] m_axi_out_13_ARSIZE;
  (* RS_HS = "m_axi_out_13_AR.valid" *)output m_axi_out_13_ARVALID;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [63:0] m_axi_out_13_AWADDR;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [1:0] m_axi_out_13_AWBURST;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [3:0] m_axi_out_13_AWCACHE;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [0:0] m_axi_out_13_AWID;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [7:0] m_axi_out_13_AWLEN;
  (* RS_HS = "m_axi_out_13_AW.data" *)output m_axi_out_13_AWLOCK;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [2:0] m_axi_out_13_AWPROT;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [3:0] m_axi_out_13_AWQOS;
  (* RS_HS = "m_axi_out_13_AW.ready" *)input m_axi_out_13_AWREADY;
  (* RS_HS = "m_axi_out_13_AW.data" *)output [2:0] m_axi_out_13_AWSIZE;
  (* RS_HS = "m_axi_out_13_AW.valid" *)output m_axi_out_13_AWVALID;
  (* RS_HS = "m_axi_out_13_B.data" *)input [0:0] m_axi_out_13_BID;
  (* RS_HS = "m_axi_out_13_B.ready" *)output m_axi_out_13_BREADY;
  (* RS_HS = "m_axi_out_13_B.data" *)input [1:0] m_axi_out_13_BRESP;
  (* RS_HS = "m_axi_out_13_B.valid" *)input m_axi_out_13_BVALID;
  (* RS_HS = "m_axi_out_13_R.data" *)input [511:0] m_axi_out_13_RDATA;
  (* RS_HS = "m_axi_out_13_R.data" *)input [0:0] m_axi_out_13_RID;
  (* RS_HS = "m_axi_out_13_R.data" *)input m_axi_out_13_RLAST;
  (* RS_HS = "m_axi_out_13_R.ready" *)output m_axi_out_13_RREADY;
  (* RS_HS = "m_axi_out_13_R.data" *)input [1:0] m_axi_out_13_RRESP;
  (* RS_HS = "m_axi_out_13_R.valid" *)input m_axi_out_13_RVALID;
  (* RS_HS = "m_axi_out_13_W.data" *)output [511:0] m_axi_out_13_WDATA;
  (* RS_HS = "m_axi_out_13_W.data" *)output m_axi_out_13_WLAST;
  (* RS_HS = "m_axi_out_13_W.ready" *)input m_axi_out_13_WREADY;
  (* RS_HS = "m_axi_out_13_W.data" *)output [63:0] m_axi_out_13_WSTRB;
  (* RS_HS = "m_axi_out_13_W.valid" *)output m_axi_out_13_WVALID;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [63:0] m_axi_in_14_ARADDR;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [1:0] m_axi_in_14_ARBURST;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [3:0] m_axi_in_14_ARCACHE;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [0:0] m_axi_in_14_ARID;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [7:0] m_axi_in_14_ARLEN;
  (* RS_HS = "m_axi_in_14_AR.data" *)output m_axi_in_14_ARLOCK;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [2:0] m_axi_in_14_ARPROT;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [3:0] m_axi_in_14_ARQOS;
  (* RS_HS = "m_axi_in_14_AR.ready" *)input m_axi_in_14_ARREADY;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [2:0] m_axi_in_14_ARSIZE;
  (* RS_HS = "m_axi_in_14_AR.valid" *)output m_axi_in_14_ARVALID;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [63:0] m_axi_in_14_AWADDR;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [1:0] m_axi_in_14_AWBURST;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [3:0] m_axi_in_14_AWCACHE;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [0:0] m_axi_in_14_AWID;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [7:0] m_axi_in_14_AWLEN;
  (* RS_HS = "m_axi_in_14_AW.data" *)output m_axi_in_14_AWLOCK;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [2:0] m_axi_in_14_AWPROT;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [3:0] m_axi_in_14_AWQOS;
  (* RS_HS = "m_axi_in_14_AW.ready" *)input m_axi_in_14_AWREADY;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [2:0] m_axi_in_14_AWSIZE;
  (* RS_HS = "m_axi_in_14_AW.valid" *)output m_axi_in_14_AWVALID;
  (* RS_HS = "m_axi_in_14_B.data" *)input [0:0] m_axi_in_14_BID;
  (* RS_HS = "m_axi_in_14_B.ready" *)output m_axi_in_14_BREADY;
  (* RS_HS = "m_axi_in_14_B.data" *)input [1:0] m_axi_in_14_BRESP;
  (* RS_HS = "m_axi_in_14_B.valid" *)input m_axi_in_14_BVALID;
  (* RS_HS = "m_axi_in_14_R.data" *)input [511:0] m_axi_in_14_RDATA;
  (* RS_HS = "m_axi_in_14_R.data" *)input [0:0] m_axi_in_14_RID;
  (* RS_HS = "m_axi_in_14_R.data" *)input m_axi_in_14_RLAST;
  (* RS_HS = "m_axi_in_14_R.ready" *)output m_axi_in_14_RREADY;
  (* RS_HS = "m_axi_in_14_R.data" *)input [1:0] m_axi_in_14_RRESP;
  (* RS_HS = "m_axi_in_14_R.valid" *)input m_axi_in_14_RVALID;
  (* RS_HS = "m_axi_in_14_W.data" *)output [511:0] m_axi_in_14_WDATA;
  (* RS_HS = "m_axi_in_14_W.data" *)output m_axi_in_14_WLAST;
  (* RS_HS = "m_axi_in_14_W.ready" *)input m_axi_in_14_WREADY;
  (* RS_HS = "m_axi_in_14_W.data" *)output [63:0] m_axi_in_14_WSTRB;
  (* RS_HS = "m_axi_in_14_W.valid" *)output m_axi_in_14_WVALID;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [63:0] m_axi_out_14_ARADDR;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [1:0] m_axi_out_14_ARBURST;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [3:0] m_axi_out_14_ARCACHE;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [0:0] m_axi_out_14_ARID;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [7:0] m_axi_out_14_ARLEN;
  (* RS_HS = "m_axi_out_14_AR.data" *)output m_axi_out_14_ARLOCK;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [2:0] m_axi_out_14_ARPROT;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [3:0] m_axi_out_14_ARQOS;
  (* RS_HS = "m_axi_out_14_AR.ready" *)input m_axi_out_14_ARREADY;
  (* RS_HS = "m_axi_out_14_AR.data" *)output [2:0] m_axi_out_14_ARSIZE;
  (* RS_HS = "m_axi_out_14_AR.valid" *)output m_axi_out_14_ARVALID;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [63:0] m_axi_out_14_AWADDR;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [1:0] m_axi_out_14_AWBURST;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [3:0] m_axi_out_14_AWCACHE;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [0:0] m_axi_out_14_AWID;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [7:0] m_axi_out_14_AWLEN;
  (* RS_HS = "m_axi_out_14_AW.data" *)output m_axi_out_14_AWLOCK;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [2:0] m_axi_out_14_AWPROT;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [3:0] m_axi_out_14_AWQOS;
  (* RS_HS = "m_axi_out_14_AW.ready" *)input m_axi_out_14_AWREADY;
  (* RS_HS = "m_axi_out_14_AW.data" *)output [2:0] m_axi_out_14_AWSIZE;
  (* RS_HS = "m_axi_out_14_AW.valid" *)output m_axi_out_14_AWVALID;
  (* RS_HS = "m_axi_out_14_B.data" *)input [0:0] m_axi_out_14_BID;
  (* RS_HS = "m_axi_out_14_B.ready" *)output m_axi_out_14_BREADY;
  (* RS_HS = "m_axi_out_14_B.data" *)input [1:0] m_axi_out_14_BRESP;
  (* RS_HS = "m_axi_out_14_B.valid" *)input m_axi_out_14_BVALID;
  (* RS_HS = "m_axi_out_14_R.data" *)input [511:0] m_axi_out_14_RDATA;
  (* RS_HS = "m_axi_out_14_R.data" *)input [0:0] m_axi_out_14_RID;
  (* RS_HS = "m_axi_out_14_R.data" *)input m_axi_out_14_RLAST;
  (* RS_HS = "m_axi_out_14_R.ready" *)output m_axi_out_14_RREADY;
  (* RS_HS = "m_axi_out_14_R.data" *)input [1:0] m_axi_out_14_RRESP;
  (* RS_HS = "m_axi_out_14_R.valid" *)input m_axi_out_14_RVALID;
  (* RS_HS = "m_axi_out_14_W.data" *)output [511:0] m_axi_out_14_WDATA;
  (* RS_HS = "m_axi_out_14_W.data" *)output m_axi_out_14_WLAST;
  (* RS_HS = "m_axi_out_14_W.ready" *)input m_axi_out_14_WREADY;
  (* RS_HS = "m_axi_out_14_W.data" *)output [63:0] m_axi_out_14_WSTRB;
  (* RS_HS = "m_axi_out_14_W.valid" *)output m_axi_out_14_WVALID;
  wire ap_start;
  wire [63:0] in_0;
  wire [63:0] out_0;
  wire [63:0] in_1;
  wire [63:0] out_1;
  wire [63:0] in_2;
  wire [63:0] out_2;
  wire [63:0] in_3;
  wire [63:0] out_3;
  wire [63:0] in_4;
  wire [63:0] out_4;
  wire [63:0] in_5;
  wire [63:0] out_5;
  wire [63:0] in_6;
  wire [63:0] out_6;
  wire [63:0] in_7;
  wire [63:0] out_7;
  wire [63:0] in_8;
  wire [63:0] out_8;
  wire [63:0] in_9;
  wire [63:0] out_9;
  wire [63:0] in_10;
  wire [63:0] out_10;
  wire [63:0] in_11;
  wire [63:0] out_11;
  wire [63:0] in_12;
  wire [63:0] out_12;
  wire [63:0] in_13;
  wire [63:0] out_13;
  wire [63:0] in_14;
  wire [63:0] out_14;
  wire [31:0] iters;
  wire [512:0] k_rd_unikernel_0__dout;
  wire k_rd_unikernel_0__empty_n;
  wire k_rd_unikernel_0__read;
  wire [512:0] k_rd_unikernel_0__din;
  wire k_rd_unikernel_0__full_n;
  wire k_rd_unikernel_0__write;
  wire [512:0] k_rd_unikernel_10__dout;
  wire k_rd_unikernel_10__empty_n;
  wire k_rd_unikernel_10__read;
  wire [512:0] k_rd_unikernel_10__din;
  wire k_rd_unikernel_10__full_n;
  wire k_rd_unikernel_10__write;
  wire [512:0] k_rd_unikernel_11__dout;
  wire k_rd_unikernel_11__empty_n;
  wire k_rd_unikernel_11__read;
  wire [512:0] k_rd_unikernel_11__din;
  wire k_rd_unikernel_11__full_n;
  wire k_rd_unikernel_11__write;
  wire [512:0] k_rd_unikernel_12__dout;
  wire k_rd_unikernel_12__empty_n;
  wire k_rd_unikernel_12__read;
  wire [512:0] k_rd_unikernel_12__din;
  wire k_rd_unikernel_12__full_n;
  wire k_rd_unikernel_12__write;
  wire [512:0] k_rd_unikernel_13__dout;
  wire k_rd_unikernel_13__empty_n;
  wire k_rd_unikernel_13__read;
  wire [512:0] k_rd_unikernel_13__din;
  wire k_rd_unikernel_13__full_n;
  wire k_rd_unikernel_13__write;
  wire [512:0] k_rd_unikernel_14__dout;
  wire k_rd_unikernel_14__empty_n;
  wire k_rd_unikernel_14__read;
  wire [512:0] k_rd_unikernel_14__din;
  wire k_rd_unikernel_14__full_n;
  wire k_rd_unikernel_14__write;
  wire [512:0] k_rd_unikernel_1__dout;
  wire k_rd_unikernel_1__empty_n;
  wire k_rd_unikernel_1__read;
  wire [512:0] k_rd_unikernel_1__din;
  wire k_rd_unikernel_1__full_n;
  wire k_rd_unikernel_1__write;
  wire [512:0] k_rd_unikernel_2__dout;
  wire k_rd_unikernel_2__empty_n;
  wire k_rd_unikernel_2__read;
  wire [512:0] k_rd_unikernel_2__din;
  wire k_rd_unikernel_2__full_n;
  wire k_rd_unikernel_2__write;
  wire [512:0] k_rd_unikernel_3__dout;
  wire k_rd_unikernel_3__empty_n;
  wire k_rd_unikernel_3__read;
  wire [512:0] k_rd_unikernel_3__din;
  wire k_rd_unikernel_3__full_n;
  wire k_rd_unikernel_3__write;
  wire [512:0] k_rd_unikernel_4__dout;
  wire k_rd_unikernel_4__empty_n;
  wire k_rd_unikernel_4__read;
  wire [512:0] k_rd_unikernel_4__din;
  wire k_rd_unikernel_4__full_n;
  wire k_rd_unikernel_4__write;
  wire [512:0] k_rd_unikernel_5__dout;
  wire k_rd_unikernel_5__empty_n;
  wire k_rd_unikernel_5__read;
  wire [512:0] k_rd_unikernel_5__din;
  wire k_rd_unikernel_5__full_n;
  wire k_rd_unikernel_5__write;
  wire [512:0] k_rd_unikernel_6__dout;
  wire k_rd_unikernel_6__empty_n;
  wire k_rd_unikernel_6__read;
  wire [512:0] k_rd_unikernel_6__din;
  wire k_rd_unikernel_6__full_n;
  wire k_rd_unikernel_6__write;
  wire [512:0] k_rd_unikernel_7__dout;
  wire k_rd_unikernel_7__empty_n;
  wire k_rd_unikernel_7__read;
  wire [512:0] k_rd_unikernel_7__din;
  wire k_rd_unikernel_7__full_n;
  wire k_rd_unikernel_7__write;
  wire [512:0] k_rd_unikernel_8__dout;
  wire k_rd_unikernel_8__empty_n;
  wire k_rd_unikernel_8__read;
  wire [512:0] k_rd_unikernel_8__din;
  wire k_rd_unikernel_8__full_n;
  wire k_rd_unikernel_8__write;
  wire [512:0] k_rd_unikernel_9__dout;
  wire k_rd_unikernel_9__empty_n;
  wire k_rd_unikernel_9__read;
  wire [512:0] k_rd_unikernel_9__din;
  wire k_rd_unikernel_9__full_n;
  wire k_rd_unikernel_9__write;
  wire [512:0] k_wr_unikernel_0__dout;
  wire k_wr_unikernel_0__empty_n;
  wire k_wr_unikernel_0__read;
  wire [512:0] k_wr_unikernel_0__din;
  wire k_wr_unikernel_0__full_n;
  wire k_wr_unikernel_0__write;
  wire [512:0] k_wr_unikernel_10__dout;
  wire k_wr_unikernel_10__empty_n;
  wire k_wr_unikernel_10__read;
  wire [512:0] k_wr_unikernel_10__din;
  wire k_wr_unikernel_10__full_n;
  wire k_wr_unikernel_10__write;
  wire [512:0] k_wr_unikernel_11__dout;
  wire k_wr_unikernel_11__empty_n;
  wire k_wr_unikernel_11__read;
  wire [512:0] k_wr_unikernel_11__din;
  wire k_wr_unikernel_11__full_n;
  wire k_wr_unikernel_11__write;
  wire [512:0] k_wr_unikernel_12__dout;
  wire k_wr_unikernel_12__empty_n;
  wire k_wr_unikernel_12__read;
  wire [512:0] k_wr_unikernel_12__din;
  wire k_wr_unikernel_12__full_n;
  wire k_wr_unikernel_12__write;
  wire [512:0] k_wr_unikernel_13__dout;
  wire k_wr_unikernel_13__empty_n;
  wire k_wr_unikernel_13__read;
  wire [512:0] k_wr_unikernel_13__din;
  wire k_wr_unikernel_13__full_n;
  wire k_wr_unikernel_13__write;
  wire [512:0] k_wr_unikernel_14__dout;
  wire k_wr_unikernel_14__empty_n;
  wire k_wr_unikernel_14__read;
  wire [512:0] k_wr_unikernel_14__din;
  wire k_wr_unikernel_14__full_n;
  wire k_wr_unikernel_14__write;
  wire [512:0] k_wr_unikernel_1__dout;
  wire k_wr_unikernel_1__empty_n;
  wire k_wr_unikernel_1__read;
  wire [512:0] k_wr_unikernel_1__din;
  wire k_wr_unikernel_1__full_n;
  wire k_wr_unikernel_1__write;
  wire [512:0] k_wr_unikernel_2__dout;
  wire k_wr_unikernel_2__empty_n;
  wire k_wr_unikernel_2__read;
  wire [512:0] k_wr_unikernel_2__din;
  wire k_wr_unikernel_2__full_n;
  wire k_wr_unikernel_2__write;
  wire [512:0] k_wr_unikernel_3__dout;
  wire k_wr_unikernel_3__empty_n;
  wire k_wr_unikernel_3__read;
  wire [512:0] k_wr_unikernel_3__din;
  wire k_wr_unikernel_3__full_n;
  wire k_wr_unikernel_3__write;
  wire [512:0] k_wr_unikernel_4__dout;
  wire k_wr_unikernel_4__empty_n;
  wire k_wr_unikernel_4__read;
  wire [512:0] k_wr_unikernel_4__din;
  wire k_wr_unikernel_4__full_n;
  wire k_wr_unikernel_4__write;
  wire [512:0] k_wr_unikernel_5__dout;
  wire k_wr_unikernel_5__empty_n;
  wire k_wr_unikernel_5__read;
  wire [512:0] k_wr_unikernel_5__din;
  wire k_wr_unikernel_5__full_n;
  wire k_wr_unikernel_5__write;
  wire [512:0] k_wr_unikernel_6__dout;
  wire k_wr_unikernel_6__empty_n;
  wire k_wr_unikernel_6__read;
  wire [512:0] k_wr_unikernel_6__din;
  wire k_wr_unikernel_6__full_n;
  wire k_wr_unikernel_6__write;
  wire [512:0] k_wr_unikernel_7__dout;
  wire k_wr_unikernel_7__empty_n;
  wire k_wr_unikernel_7__read;
  wire [512:0] k_wr_unikernel_7__din;
  wire k_wr_unikernel_7__full_n;
  wire k_wr_unikernel_7__write;
  wire [512:0] k_wr_unikernel_8__dout;
  wire k_wr_unikernel_8__empty_n;
  wire k_wr_unikernel_8__read;
  wire [512:0] k_wr_unikernel_8__din;
  wire k_wr_unikernel_8__full_n;
  wire k_wr_unikernel_8__write;
  wire [512:0] k_wr_unikernel_9__dout;
  wire k_wr_unikernel_9__empty_n;
  wire k_wr_unikernel_9__read;
  wire [512:0] k_wr_unikernel_9__din;
  wire k_wr_unikernel_9__full_n;
  wire k_wr_unikernel_9__write;
  wire [31:0] JACOBI3D_0___iters__q0;
  wire JACOBI3D_0__ap_start;
  wire JACOBI3D_0__ap_ready;
  wire JACOBI3D_0__ap_done;
  wire JACOBI3D_0__ap_idle;
  wire [31:0] JACOBI3D_1___iters__q0;
  wire JACOBI3D_1__ap_start;
  wire JACOBI3D_1__ap_ready;
  wire JACOBI3D_1__ap_done;
  wire JACOBI3D_1__ap_idle;
  wire [31:0] JACOBI3D_2___iters__q0;
  wire JACOBI3D_2__ap_start;
  wire JACOBI3D_2__ap_ready;
  wire JACOBI3D_2__ap_done;
  wire JACOBI3D_2__ap_idle;
  wire [31:0] JACOBI3D_3___iters__q0;
  wire JACOBI3D_3__ap_start;
  wire JACOBI3D_3__ap_ready;
  wire JACOBI3D_3__ap_done;
  wire JACOBI3D_3__ap_idle;
  wire [31:0] JACOBI3D_4___iters__q0;
  wire JACOBI3D_4__ap_start;
  wire JACOBI3D_4__ap_ready;
  wire JACOBI3D_4__ap_done;
  wire JACOBI3D_4__ap_idle;
  wire [31:0] JACOBI3D_5___iters__q0;
  wire JACOBI3D_5__ap_start;
  wire JACOBI3D_5__ap_ready;
  wire JACOBI3D_5__ap_done;
  wire JACOBI3D_5__ap_idle;
  wire [31:0] JACOBI3D_6___iters__q0;
  wire JACOBI3D_6__ap_start;
  wire JACOBI3D_6__ap_ready;
  wire JACOBI3D_6__ap_done;
  wire JACOBI3D_6__ap_idle;
  wire [31:0] JACOBI3D_7___iters__q0;
  wire JACOBI3D_7__ap_start;
  wire JACOBI3D_7__ap_ready;
  wire JACOBI3D_7__ap_done;
  wire JACOBI3D_7__ap_idle;
  wire [31:0] JACOBI3D_8___iters__q0;
  wire JACOBI3D_8__ap_start;
  wire JACOBI3D_8__ap_ready;
  wire JACOBI3D_8__ap_done;
  wire JACOBI3D_8__ap_idle;
  wire [31:0] JACOBI3D_9___iters__q0;
  wire JACOBI3D_9__ap_start;
  wire JACOBI3D_9__ap_ready;
  wire JACOBI3D_9__ap_done;
  wire JACOBI3D_9__ap_idle;
  wire [31:0] JACOBI3D_10___iters__q0;
  wire JACOBI3D_10__ap_start;
  wire JACOBI3D_10__ap_ready;
  wire JACOBI3D_10__ap_done;
  wire JACOBI3D_10__ap_idle;
  wire [31:0] JACOBI3D_11___iters__q0;
  wire JACOBI3D_11__ap_start;
  wire JACOBI3D_11__ap_ready;
  wire JACOBI3D_11__ap_done;
  wire JACOBI3D_11__ap_idle;
  wire [31:0] JACOBI3D_12___iters__q0;
  wire JACOBI3D_12__ap_start;
  wire JACOBI3D_12__ap_ready;
  wire JACOBI3D_12__ap_done;
  wire JACOBI3D_12__ap_idle;
  wire [31:0] JACOBI3D_13___iters__q0;
  wire JACOBI3D_13__ap_start;
  wire JACOBI3D_13__ap_ready;
  wire JACOBI3D_13__ap_done;
  wire JACOBI3D_13__ap_idle;
  wire [31:0] JACOBI3D_14___iters__q0;
  wire JACOBI3D_14__ap_start;
  wire JACOBI3D_14__ap_ready;
  wire JACOBI3D_14__ap_done;
  wire JACOBI3D_14__ap_idle;
  wire [63:0] inter_kernel_0___in_0__q0;
  wire [63:0] in_0_read_addr__din;
  wire in_0_read_addr__full_n;
  wire in_0_read_addr__write;
  wire [511:0] in_0_read_data__dout;
  wire in_0_read_data__empty_n;
  wire in_0_read_data__read;
  wire [63:0] in_0_write_addr__din;
  wire in_0_write_addr__full_n;
  wire in_0_write_addr__write;
  wire [511:0] in_0_write_data__din;
  wire in_0_write_data__full_n;
  wire in_0_write_data__write;
  wire [7:0] in_0_write_resp__dout;
  wire in_0_write_resp__empty_n;
  wire in_0_write_resp__read;
  wire [31:0] inter_kernel_0___iters__q0;
  wire [63:0] inter_kernel_0___out_0__q0;
  wire [63:0] out_0_read_addr__din;
  wire out_0_read_addr__full_n;
  wire out_0_read_addr__write;
  wire [511:0] out_0_read_data__dout;
  wire out_0_read_data__empty_n;
  wire out_0_read_data__read;
  wire [63:0] out_0_write_addr__din;
  wire out_0_write_addr__full_n;
  wire out_0_write_addr__write;
  wire [511:0] out_0_write_data__din;
  wire out_0_write_data__full_n;
  wire out_0_write_data__write;
  wire [7:0] out_0_write_resp__dout;
  wire out_0_write_resp__empty_n;
  wire out_0_write_resp__read;
  wire inter_kernel_0__ap_start;
  wire inter_kernel_0__ap_ready;
  wire inter_kernel_0__ap_done;
  wire inter_kernel_0__ap_idle;
  wire [63:0] inter_kernel_1___in_1__q0;
  wire [63:0] in_1_read_addr__din;
  wire in_1_read_addr__full_n;
  wire in_1_read_addr__write;
  wire [511:0] in_1_read_data__dout;
  wire in_1_read_data__empty_n;
  wire in_1_read_data__read;
  wire [63:0] in_1_write_addr__din;
  wire in_1_write_addr__full_n;
  wire in_1_write_addr__write;
  wire [511:0] in_1_write_data__din;
  wire in_1_write_data__full_n;
  wire in_1_write_data__write;
  wire [7:0] in_1_write_resp__dout;
  wire in_1_write_resp__empty_n;
  wire in_1_write_resp__read;
  wire [31:0] inter_kernel_1___iters__q0;
  wire [63:0] inter_kernel_1___out_1__q0;
  wire [63:0] out_1_read_addr__din;
  wire out_1_read_addr__full_n;
  wire out_1_read_addr__write;
  wire [511:0] out_1_read_data__dout;
  wire out_1_read_data__empty_n;
  wire out_1_read_data__read;
  wire [63:0] out_1_write_addr__din;
  wire out_1_write_addr__full_n;
  wire out_1_write_addr__write;
  wire [511:0] out_1_write_data__din;
  wire out_1_write_data__full_n;
  wire out_1_write_data__write;
  wire [7:0] out_1_write_resp__dout;
  wire out_1_write_resp__empty_n;
  wire out_1_write_resp__read;
  wire inter_kernel_1__ap_start;
  wire inter_kernel_1__ap_ready;
  wire inter_kernel_1__ap_done;
  wire inter_kernel_1__ap_idle;
  wire [63:0] inter_kernel_2___in_2__q0;
  wire [63:0] in_2_read_addr__din;
  wire in_2_read_addr__full_n;
  wire in_2_read_addr__write;
  wire [511:0] in_2_read_data__dout;
  wire in_2_read_data__empty_n;
  wire in_2_read_data__read;
  wire [63:0] in_2_write_addr__din;
  wire in_2_write_addr__full_n;
  wire in_2_write_addr__write;
  wire [511:0] in_2_write_data__din;
  wire in_2_write_data__full_n;
  wire in_2_write_data__write;
  wire [7:0] in_2_write_resp__dout;
  wire in_2_write_resp__empty_n;
  wire in_2_write_resp__read;
  wire [31:0] inter_kernel_2___iters__q0;
  wire [63:0] inter_kernel_2___out_2__q0;
  wire [63:0] out_2_read_addr__din;
  wire out_2_read_addr__full_n;
  wire out_2_read_addr__write;
  wire [511:0] out_2_read_data__dout;
  wire out_2_read_data__empty_n;
  wire out_2_read_data__read;
  wire [63:0] out_2_write_addr__din;
  wire out_2_write_addr__full_n;
  wire out_2_write_addr__write;
  wire [511:0] out_2_write_data__din;
  wire out_2_write_data__full_n;
  wire out_2_write_data__write;
  wire [7:0] out_2_write_resp__dout;
  wire out_2_write_resp__empty_n;
  wire out_2_write_resp__read;
  wire inter_kernel_2__ap_start;
  wire inter_kernel_2__ap_ready;
  wire inter_kernel_2__ap_done;
  wire inter_kernel_2__ap_idle;
  wire [63:0] inter_kernel_3___in_3__q0;
  wire [63:0] in_3_read_addr__din;
  wire in_3_read_addr__full_n;
  wire in_3_read_addr__write;
  wire [511:0] in_3_read_data__dout;
  wire in_3_read_data__empty_n;
  wire in_3_read_data__read;
  wire [63:0] in_3_write_addr__din;
  wire in_3_write_addr__full_n;
  wire in_3_write_addr__write;
  wire [511:0] in_3_write_data__din;
  wire in_3_write_data__full_n;
  wire in_3_write_data__write;
  wire [7:0] in_3_write_resp__dout;
  wire in_3_write_resp__empty_n;
  wire in_3_write_resp__read;
  wire [31:0] inter_kernel_3___iters__q0;
  wire [63:0] inter_kernel_3___out_3__q0;
  wire [63:0] out_3_read_addr__din;
  wire out_3_read_addr__full_n;
  wire out_3_read_addr__write;
  wire [511:0] out_3_read_data__dout;
  wire out_3_read_data__empty_n;
  wire out_3_read_data__read;
  wire [63:0] out_3_write_addr__din;
  wire out_3_write_addr__full_n;
  wire out_3_write_addr__write;
  wire [511:0] out_3_write_data__din;
  wire out_3_write_data__full_n;
  wire out_3_write_data__write;
  wire [7:0] out_3_write_resp__dout;
  wire out_3_write_resp__empty_n;
  wire out_3_write_resp__read;
  wire inter_kernel_3__ap_start;
  wire inter_kernel_3__ap_ready;
  wire inter_kernel_3__ap_done;
  wire inter_kernel_3__ap_idle;
  wire [63:0] inter_kernel_4___in_4__q0;
  wire [63:0] in_4_read_addr__din;
  wire in_4_read_addr__full_n;
  wire in_4_read_addr__write;
  wire [511:0] in_4_read_data__dout;
  wire in_4_read_data__empty_n;
  wire in_4_read_data__read;
  wire [63:0] in_4_write_addr__din;
  wire in_4_write_addr__full_n;
  wire in_4_write_addr__write;
  wire [511:0] in_4_write_data__din;
  wire in_4_write_data__full_n;
  wire in_4_write_data__write;
  wire [7:0] in_4_write_resp__dout;
  wire in_4_write_resp__empty_n;
  wire in_4_write_resp__read;
  wire [31:0] inter_kernel_4___iters__q0;
  wire [63:0] inter_kernel_4___out_4__q0;
  wire [63:0] out_4_read_addr__din;
  wire out_4_read_addr__full_n;
  wire out_4_read_addr__write;
  wire [511:0] out_4_read_data__dout;
  wire out_4_read_data__empty_n;
  wire out_4_read_data__read;
  wire [63:0] out_4_write_addr__din;
  wire out_4_write_addr__full_n;
  wire out_4_write_addr__write;
  wire [511:0] out_4_write_data__din;
  wire out_4_write_data__full_n;
  wire out_4_write_data__write;
  wire [7:0] out_4_write_resp__dout;
  wire out_4_write_resp__empty_n;
  wire out_4_write_resp__read;
  wire inter_kernel_4__ap_start;
  wire inter_kernel_4__ap_ready;
  wire inter_kernel_4__ap_done;
  wire inter_kernel_4__ap_idle;
  wire [63:0] inter_kernel_5___in_5__q0;
  wire [63:0] in_5_read_addr__din;
  wire in_5_read_addr__full_n;
  wire in_5_read_addr__write;
  wire [511:0] in_5_read_data__dout;
  wire in_5_read_data__empty_n;
  wire in_5_read_data__read;
  wire [63:0] in_5_write_addr__din;
  wire in_5_write_addr__full_n;
  wire in_5_write_addr__write;
  wire [511:0] in_5_write_data__din;
  wire in_5_write_data__full_n;
  wire in_5_write_data__write;
  wire [7:0] in_5_write_resp__dout;
  wire in_5_write_resp__empty_n;
  wire in_5_write_resp__read;
  wire [31:0] inter_kernel_5___iters__q0;
  wire [63:0] inter_kernel_5___out_5__q0;
  wire [63:0] out_5_read_addr__din;
  wire out_5_read_addr__full_n;
  wire out_5_read_addr__write;
  wire [511:0] out_5_read_data__dout;
  wire out_5_read_data__empty_n;
  wire out_5_read_data__read;
  wire [63:0] out_5_write_addr__din;
  wire out_5_write_addr__full_n;
  wire out_5_write_addr__write;
  wire [511:0] out_5_write_data__din;
  wire out_5_write_data__full_n;
  wire out_5_write_data__write;
  wire [7:0] out_5_write_resp__dout;
  wire out_5_write_resp__empty_n;
  wire out_5_write_resp__read;
  wire inter_kernel_5__ap_start;
  wire inter_kernel_5__ap_ready;
  wire inter_kernel_5__ap_done;
  wire inter_kernel_5__ap_idle;
  wire [63:0] inter_kernel_6___in_6__q0;
  wire [63:0] in_6_read_addr__din;
  wire in_6_read_addr__full_n;
  wire in_6_read_addr__write;
  wire [511:0] in_6_read_data__dout;
  wire in_6_read_data__empty_n;
  wire in_6_read_data__read;
  wire [63:0] in_6_write_addr__din;
  wire in_6_write_addr__full_n;
  wire in_6_write_addr__write;
  wire [511:0] in_6_write_data__din;
  wire in_6_write_data__full_n;
  wire in_6_write_data__write;
  wire [7:0] in_6_write_resp__dout;
  wire in_6_write_resp__empty_n;
  wire in_6_write_resp__read;
  wire [31:0] inter_kernel_6___iters__q0;
  wire [63:0] inter_kernel_6___out_6__q0;
  wire [63:0] out_6_read_addr__din;
  wire out_6_read_addr__full_n;
  wire out_6_read_addr__write;
  wire [511:0] out_6_read_data__dout;
  wire out_6_read_data__empty_n;
  wire out_6_read_data__read;
  wire [63:0] out_6_write_addr__din;
  wire out_6_write_addr__full_n;
  wire out_6_write_addr__write;
  wire [511:0] out_6_write_data__din;
  wire out_6_write_data__full_n;
  wire out_6_write_data__write;
  wire [7:0] out_6_write_resp__dout;
  wire out_6_write_resp__empty_n;
  wire out_6_write_resp__read;
  wire inter_kernel_6__ap_start;
  wire inter_kernel_6__ap_ready;
  wire inter_kernel_6__ap_done;
  wire inter_kernel_6__ap_idle;
  wire [63:0] inter_kernel_7___in_7__q0;
  wire [63:0] in_7_read_addr__din;
  wire in_7_read_addr__full_n;
  wire in_7_read_addr__write;
  wire [511:0] in_7_read_data__dout;
  wire in_7_read_data__empty_n;
  wire in_7_read_data__read;
  wire [63:0] in_7_write_addr__din;
  wire in_7_write_addr__full_n;
  wire in_7_write_addr__write;
  wire [511:0] in_7_write_data__din;
  wire in_7_write_data__full_n;
  wire in_7_write_data__write;
  wire [7:0] in_7_write_resp__dout;
  wire in_7_write_resp__empty_n;
  wire in_7_write_resp__read;
  wire [31:0] inter_kernel_7___iters__q0;
  wire [63:0] inter_kernel_7___out_7__q0;
  wire [63:0] out_7_read_addr__din;
  wire out_7_read_addr__full_n;
  wire out_7_read_addr__write;
  wire [511:0] out_7_read_data__dout;
  wire out_7_read_data__empty_n;
  wire out_7_read_data__read;
  wire [63:0] out_7_write_addr__din;
  wire out_7_write_addr__full_n;
  wire out_7_write_addr__write;
  wire [511:0] out_7_write_data__din;
  wire out_7_write_data__full_n;
  wire out_7_write_data__write;
  wire [7:0] out_7_write_resp__dout;
  wire out_7_write_resp__empty_n;
  wire out_7_write_resp__read;
  wire inter_kernel_7__ap_start;
  wire inter_kernel_7__ap_ready;
  wire inter_kernel_7__ap_done;
  wire inter_kernel_7__ap_idle;
  wire [63:0] inter_kernel_8___in_8__q0;
  wire [63:0] in_8_read_addr__din;
  wire in_8_read_addr__full_n;
  wire in_8_read_addr__write;
  wire [511:0] in_8_read_data__dout;
  wire in_8_read_data__empty_n;
  wire in_8_read_data__read;
  wire [63:0] in_8_write_addr__din;
  wire in_8_write_addr__full_n;
  wire in_8_write_addr__write;
  wire [511:0] in_8_write_data__din;
  wire in_8_write_data__full_n;
  wire in_8_write_data__write;
  wire [7:0] in_8_write_resp__dout;
  wire in_8_write_resp__empty_n;
  wire in_8_write_resp__read;
  wire [31:0] inter_kernel_8___iters__q0;
  wire [63:0] inter_kernel_8___out_8__q0;
  wire [63:0] out_8_read_addr__din;
  wire out_8_read_addr__full_n;
  wire out_8_read_addr__write;
  wire [511:0] out_8_read_data__dout;
  wire out_8_read_data__empty_n;
  wire out_8_read_data__read;
  wire [63:0] out_8_write_addr__din;
  wire out_8_write_addr__full_n;
  wire out_8_write_addr__write;
  wire [511:0] out_8_write_data__din;
  wire out_8_write_data__full_n;
  wire out_8_write_data__write;
  wire [7:0] out_8_write_resp__dout;
  wire out_8_write_resp__empty_n;
  wire out_8_write_resp__read;
  wire inter_kernel_8__ap_start;
  wire inter_kernel_8__ap_ready;
  wire inter_kernel_8__ap_done;
  wire inter_kernel_8__ap_idle;
  wire [63:0] inter_kernel_9___in_9__q0;
  wire [63:0] in_9_read_addr__din;
  wire in_9_read_addr__full_n;
  wire in_9_read_addr__write;
  wire [511:0] in_9_read_data__dout;
  wire in_9_read_data__empty_n;
  wire in_9_read_data__read;
  wire [63:0] in_9_write_addr__din;
  wire in_9_write_addr__full_n;
  wire in_9_write_addr__write;
  wire [511:0] in_9_write_data__din;
  wire in_9_write_data__full_n;
  wire in_9_write_data__write;
  wire [7:0] in_9_write_resp__dout;
  wire in_9_write_resp__empty_n;
  wire in_9_write_resp__read;
  wire [31:0] inter_kernel_9___iters__q0;
  wire [63:0] inter_kernel_9___out_9__q0;
  wire [63:0] out_9_read_addr__din;
  wire out_9_read_addr__full_n;
  wire out_9_read_addr__write;
  wire [511:0] out_9_read_data__dout;
  wire out_9_read_data__empty_n;
  wire out_9_read_data__read;
  wire [63:0] out_9_write_addr__din;
  wire out_9_write_addr__full_n;
  wire out_9_write_addr__write;
  wire [511:0] out_9_write_data__din;
  wire out_9_write_data__full_n;
  wire out_9_write_data__write;
  wire [7:0] out_9_write_resp__dout;
  wire out_9_write_resp__empty_n;
  wire out_9_write_resp__read;
  wire inter_kernel_9__ap_start;
  wire inter_kernel_9__ap_ready;
  wire inter_kernel_9__ap_done;
  wire inter_kernel_9__ap_idle;
  wire [63:0] inter_kernel_10___in_10__q0;
  wire [63:0] in_10_read_addr__din;
  wire in_10_read_addr__full_n;
  wire in_10_read_addr__write;
  wire [511:0] in_10_read_data__dout;
  wire in_10_read_data__empty_n;
  wire in_10_read_data__read;
  wire [63:0] in_10_write_addr__din;
  wire in_10_write_addr__full_n;
  wire in_10_write_addr__write;
  wire [511:0] in_10_write_data__din;
  wire in_10_write_data__full_n;
  wire in_10_write_data__write;
  wire [7:0] in_10_write_resp__dout;
  wire in_10_write_resp__empty_n;
  wire in_10_write_resp__read;
  wire [31:0] inter_kernel_10___iters__q0;
  wire [63:0] inter_kernel_10___out_10__q0;
  wire [63:0] out_10_read_addr__din;
  wire out_10_read_addr__full_n;
  wire out_10_read_addr__write;
  wire [511:0] out_10_read_data__dout;
  wire out_10_read_data__empty_n;
  wire out_10_read_data__read;
  wire [63:0] out_10_write_addr__din;
  wire out_10_write_addr__full_n;
  wire out_10_write_addr__write;
  wire [511:0] out_10_write_data__din;
  wire out_10_write_data__full_n;
  wire out_10_write_data__write;
  wire [7:0] out_10_write_resp__dout;
  wire out_10_write_resp__empty_n;
  wire out_10_write_resp__read;
  wire inter_kernel_10__ap_start;
  wire inter_kernel_10__ap_ready;
  wire inter_kernel_10__ap_done;
  wire inter_kernel_10__ap_idle;
  wire [63:0] inter_kernel_11___in_11__q0;
  wire [63:0] in_11_read_addr__din;
  wire in_11_read_addr__full_n;
  wire in_11_read_addr__write;
  wire [511:0] in_11_read_data__dout;
  wire in_11_read_data__empty_n;
  wire in_11_read_data__read;
  wire [63:0] in_11_write_addr__din;
  wire in_11_write_addr__full_n;
  wire in_11_write_addr__write;
  wire [511:0] in_11_write_data__din;
  wire in_11_write_data__full_n;
  wire in_11_write_data__write;
  wire [7:0] in_11_write_resp__dout;
  wire in_11_write_resp__empty_n;
  wire in_11_write_resp__read;
  wire [31:0] inter_kernel_11___iters__q0;
  wire [63:0] inter_kernel_11___out_11__q0;
  wire [63:0] out_11_read_addr__din;
  wire out_11_read_addr__full_n;
  wire out_11_read_addr__write;
  wire [511:0] out_11_read_data__dout;
  wire out_11_read_data__empty_n;
  wire out_11_read_data__read;
  wire [63:0] out_11_write_addr__din;
  wire out_11_write_addr__full_n;
  wire out_11_write_addr__write;
  wire [511:0] out_11_write_data__din;
  wire out_11_write_data__full_n;
  wire out_11_write_data__write;
  wire [7:0] out_11_write_resp__dout;
  wire out_11_write_resp__empty_n;
  wire out_11_write_resp__read;
  wire inter_kernel_11__ap_start;
  wire inter_kernel_11__ap_ready;
  wire inter_kernel_11__ap_done;
  wire inter_kernel_11__ap_idle;
  wire [63:0] inter_kernel_12___in_12__q0;
  wire [63:0] in_12_read_addr__din;
  wire in_12_read_addr__full_n;
  wire in_12_read_addr__write;
  wire [511:0] in_12_read_data__dout;
  wire in_12_read_data__empty_n;
  wire in_12_read_data__read;
  wire [63:0] in_12_write_addr__din;
  wire in_12_write_addr__full_n;
  wire in_12_write_addr__write;
  wire [511:0] in_12_write_data__din;
  wire in_12_write_data__full_n;
  wire in_12_write_data__write;
  wire [7:0] in_12_write_resp__dout;
  wire in_12_write_resp__empty_n;
  wire in_12_write_resp__read;
  wire [31:0] inter_kernel_12___iters__q0;
  wire [63:0] inter_kernel_12___out_12__q0;
  wire [63:0] out_12_read_addr__din;
  wire out_12_read_addr__full_n;
  wire out_12_read_addr__write;
  wire [511:0] out_12_read_data__dout;
  wire out_12_read_data__empty_n;
  wire out_12_read_data__read;
  wire [63:0] out_12_write_addr__din;
  wire out_12_write_addr__full_n;
  wire out_12_write_addr__write;
  wire [511:0] out_12_write_data__din;
  wire out_12_write_data__full_n;
  wire out_12_write_data__write;
  wire [7:0] out_12_write_resp__dout;
  wire out_12_write_resp__empty_n;
  wire out_12_write_resp__read;
  wire inter_kernel_12__ap_start;
  wire inter_kernel_12__ap_ready;
  wire inter_kernel_12__ap_done;
  wire inter_kernel_12__ap_idle;
  wire [63:0] inter_kernel_13___in_13__q0;
  wire [63:0] in_13_read_addr__din;
  wire in_13_read_addr__full_n;
  wire in_13_read_addr__write;
  wire [511:0] in_13_read_data__dout;
  wire in_13_read_data__empty_n;
  wire in_13_read_data__read;
  wire [63:0] in_13_write_addr__din;
  wire in_13_write_addr__full_n;
  wire in_13_write_addr__write;
  wire [511:0] in_13_write_data__din;
  wire in_13_write_data__full_n;
  wire in_13_write_data__write;
  wire [7:0] in_13_write_resp__dout;
  wire in_13_write_resp__empty_n;
  wire in_13_write_resp__read;
  wire [31:0] inter_kernel_13___iters__q0;
  wire [63:0] inter_kernel_13___out_13__q0;
  wire [63:0] out_13_read_addr__din;
  wire out_13_read_addr__full_n;
  wire out_13_read_addr__write;
  wire [511:0] out_13_read_data__dout;
  wire out_13_read_data__empty_n;
  wire out_13_read_data__read;
  wire [63:0] out_13_write_addr__din;
  wire out_13_write_addr__full_n;
  wire out_13_write_addr__write;
  wire [511:0] out_13_write_data__din;
  wire out_13_write_data__full_n;
  wire out_13_write_data__write;
  wire [7:0] out_13_write_resp__dout;
  wire out_13_write_resp__empty_n;
  wire out_13_write_resp__read;
  wire inter_kernel_13__ap_start;
  wire inter_kernel_13__ap_ready;
  wire inter_kernel_13__ap_done;
  wire inter_kernel_13__ap_idle;
  wire [63:0] inter_kernel_14___in_14__q0;
  wire [63:0] in_14_read_addr__din;
  wire in_14_read_addr__full_n;
  wire in_14_read_addr__write;
  wire [511:0] in_14_read_data__dout;
  wire in_14_read_data__empty_n;
  wire in_14_read_data__read;
  wire [63:0] in_14_write_addr__din;
  wire in_14_write_addr__full_n;
  wire in_14_write_addr__write;
  wire [511:0] in_14_write_data__din;
  wire in_14_write_data__full_n;
  wire in_14_write_data__write;
  wire [7:0] in_14_write_resp__dout;
  wire in_14_write_resp__empty_n;
  wire in_14_write_resp__read;
  wire [31:0] inter_kernel_14___iters__q0;
  wire [63:0] inter_kernel_14___out_14__q0;
  wire [63:0] out_14_read_addr__din;
  wire out_14_read_addr__full_n;
  wire out_14_read_addr__write;
  wire [511:0] out_14_read_data__dout;
  wire out_14_read_data__empty_n;
  wire out_14_read_data__read;
  wire [63:0] out_14_write_addr__din;
  wire out_14_write_addr__full_n;
  wire out_14_write_addr__write;
  wire [511:0] out_14_write_data__din;
  wire out_14_write_data__full_n;
  wire out_14_write_data__write;
  wire [7:0] out_14_write_resp__dout;
  wire out_14_write_resp__empty_n;
  wire out_14_write_resp__read;
  wire inter_kernel_14__ap_start;
  wire inter_kernel_14__ap_ready;
  wire inter_kernel_14__ap_done;
  wire inter_kernel_14__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;

  unikernel_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .in_0(in_0),
    .out_0(out_0),
    .in_1(in_1),
    .out_1(out_1),
    .in_2(in_2),
    .out_2(out_2),
    .in_3(in_3),
    .out_3(out_3),
    .in_4(in_4),
    .out_4(out_4),
    .in_5(in_5),
    .out_5(out_5),
    .in_6(in_6),
    .out_6(out_6),
    .in_7(in_7),
    .out_7(out_7),
    .in_8(in_8),
    .out_8(out_8),
    .in_9(in_9),
    .out_9(out_9),
    .in_10(in_10),
    .out_10(out_10),
    .in_11(in_11),
    .out_11(out_11),
    .in_12(in_12),
    .out_12(out_12),
    .in_13(in_13),
    .out_13(out_13),
    .in_14(in_14),
    .out_14(out_14),
    .iters(iters),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_0__dout),
    .if_empty_n(k_rd_unikernel_0__empty_n),
    .if_read(k_rd_unikernel_0__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_0__din),
    .if_full_n(k_rd_unikernel_0__full_n),
    .if_write(k_rd_unikernel_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_10__dout),
    .if_empty_n(k_rd_unikernel_10__empty_n),
    .if_read(k_rd_unikernel_10__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_10__din),
    .if_full_n(k_rd_unikernel_10__full_n),
    .if_write(k_rd_unikernel_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_11__dout),
    .if_empty_n(k_rd_unikernel_11__empty_n),
    .if_read(k_rd_unikernel_11__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_11__din),
    .if_full_n(k_rd_unikernel_11__full_n),
    .if_write(k_rd_unikernel_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_12__dout),
    .if_empty_n(k_rd_unikernel_12__empty_n),
    .if_read(k_rd_unikernel_12__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_12__din),
    .if_full_n(k_rd_unikernel_12__full_n),
    .if_write(k_rd_unikernel_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_13__dout),
    .if_empty_n(k_rd_unikernel_13__empty_n),
    .if_read(k_rd_unikernel_13__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_13__din),
    .if_full_n(k_rd_unikernel_13__full_n),
    .if_write(k_rd_unikernel_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_14__dout),
    .if_empty_n(k_rd_unikernel_14__empty_n),
    .if_read(k_rd_unikernel_14__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_14__din),
    .if_full_n(k_rd_unikernel_14__full_n),
    .if_write(k_rd_unikernel_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_1__dout),
    .if_empty_n(k_rd_unikernel_1__empty_n),
    .if_read(k_rd_unikernel_1__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_1__din),
    .if_full_n(k_rd_unikernel_1__full_n),
    .if_write(k_rd_unikernel_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_2__dout),
    .if_empty_n(k_rd_unikernel_2__empty_n),
    .if_read(k_rd_unikernel_2__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_2__din),
    .if_full_n(k_rd_unikernel_2__full_n),
    .if_write(k_rd_unikernel_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_3__dout),
    .if_empty_n(k_rd_unikernel_3__empty_n),
    .if_read(k_rd_unikernel_3__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_3__din),
    .if_full_n(k_rd_unikernel_3__full_n),
    .if_write(k_rd_unikernel_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_4__dout),
    .if_empty_n(k_rd_unikernel_4__empty_n),
    .if_read(k_rd_unikernel_4__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_4__din),
    .if_full_n(k_rd_unikernel_4__full_n),
    .if_write(k_rd_unikernel_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_5__dout),
    .if_empty_n(k_rd_unikernel_5__empty_n),
    .if_read(k_rd_unikernel_5__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_5__din),
    .if_full_n(k_rd_unikernel_5__full_n),
    .if_write(k_rd_unikernel_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_6__dout),
    .if_empty_n(k_rd_unikernel_6__empty_n),
    .if_read(k_rd_unikernel_6__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_6__din),
    .if_full_n(k_rd_unikernel_6__full_n),
    .if_write(k_rd_unikernel_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_7__dout),
    .if_empty_n(k_rd_unikernel_7__empty_n),
    .if_read(k_rd_unikernel_7__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_7__din),
    .if_full_n(k_rd_unikernel_7__full_n),
    .if_write(k_rd_unikernel_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_8__dout),
    .if_empty_n(k_rd_unikernel_8__empty_n),
    .if_read(k_rd_unikernel_8__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_8__din),
    .if_full_n(k_rd_unikernel_8__full_n),
    .if_write(k_rd_unikernel_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_rd_unikernel_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_rd_unikernel_9__dout),
    .if_empty_n(k_rd_unikernel_9__empty_n),
    .if_read(k_rd_unikernel_9__read),
    .if_read_ce(1'b1),
    .if_din(k_rd_unikernel_9__din),
    .if_full_n(k_rd_unikernel_9__full_n),
    .if_write(k_rd_unikernel_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_0__dout),
    .if_empty_n(k_wr_unikernel_0__empty_n),
    .if_read(k_wr_unikernel_0__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_0__din),
    .if_full_n(k_wr_unikernel_0__full_n),
    .if_write(k_wr_unikernel_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_10__dout),
    .if_empty_n(k_wr_unikernel_10__empty_n),
    .if_read(k_wr_unikernel_10__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_10__din),
    .if_full_n(k_wr_unikernel_10__full_n),
    .if_write(k_wr_unikernel_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_11__dout),
    .if_empty_n(k_wr_unikernel_11__empty_n),
    .if_read(k_wr_unikernel_11__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_11__din),
    .if_full_n(k_wr_unikernel_11__full_n),
    .if_write(k_wr_unikernel_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_12__dout),
    .if_empty_n(k_wr_unikernel_12__empty_n),
    .if_read(k_wr_unikernel_12__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_12__din),
    .if_full_n(k_wr_unikernel_12__full_n),
    .if_write(k_wr_unikernel_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_13__dout),
    .if_empty_n(k_wr_unikernel_13__empty_n),
    .if_read(k_wr_unikernel_13__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_13__din),
    .if_full_n(k_wr_unikernel_13__full_n),
    .if_write(k_wr_unikernel_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_14__dout),
    .if_empty_n(k_wr_unikernel_14__empty_n),
    .if_read(k_wr_unikernel_14__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_14__din),
    .if_full_n(k_wr_unikernel_14__full_n),
    .if_write(k_wr_unikernel_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_1__dout),
    .if_empty_n(k_wr_unikernel_1__empty_n),
    .if_read(k_wr_unikernel_1__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_1__din),
    .if_full_n(k_wr_unikernel_1__full_n),
    .if_write(k_wr_unikernel_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_2__dout),
    .if_empty_n(k_wr_unikernel_2__empty_n),
    .if_read(k_wr_unikernel_2__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_2__din),
    .if_full_n(k_wr_unikernel_2__full_n),
    .if_write(k_wr_unikernel_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_3__dout),
    .if_empty_n(k_wr_unikernel_3__empty_n),
    .if_read(k_wr_unikernel_3__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_3__din),
    .if_full_n(k_wr_unikernel_3__full_n),
    .if_write(k_wr_unikernel_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_4__dout),
    .if_empty_n(k_wr_unikernel_4__empty_n),
    .if_read(k_wr_unikernel_4__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_4__din),
    .if_full_n(k_wr_unikernel_4__full_n),
    .if_write(k_wr_unikernel_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_5__dout),
    .if_empty_n(k_wr_unikernel_5__empty_n),
    .if_read(k_wr_unikernel_5__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_5__din),
    .if_full_n(k_wr_unikernel_5__full_n),
    .if_write(k_wr_unikernel_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_6__dout),
    .if_empty_n(k_wr_unikernel_6__empty_n),
    .if_read(k_wr_unikernel_6__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_6__din),
    .if_full_n(k_wr_unikernel_6__full_n),
    .if_write(k_wr_unikernel_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_7__dout),
    .if_empty_n(k_wr_unikernel_7__empty_n),
    .if_read(k_wr_unikernel_7__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_7__din),
    .if_full_n(k_wr_unikernel_7__full_n),
    .if_write(k_wr_unikernel_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_8__dout),
    .if_empty_n(k_wr_unikernel_8__empty_n),
    .if_read(k_wr_unikernel_8__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_8__din),
    .if_full_n(k_wr_unikernel_8__full_n),
    .if_write(k_wr_unikernel_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(2),
    .DEPTH(3)
  )
  k_wr_unikernel_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(k_wr_unikernel_9__dout),
    .if_empty_n(k_wr_unikernel_9__empty_n),
    .if_read(k_wr_unikernel_9__read),
    .if_read_ce(1'b1),
    .if_din(k_wr_unikernel_9__din),
    .if_full_n(k_wr_unikernel_9__full_n),
    .if_write(k_wr_unikernel_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_0__ap_start),
    .ap_done(JACOBI3D_0__ap_done),
    .ap_idle(JACOBI3D_0__ap_idle),
    .ap_ready(JACOBI3D_0__ap_ready),
    .iters(JACOBI3D_0___iters__q0),
    .t1_s_dout(k_rd_unikernel_0__dout),
    .t1_peek_dout(k_rd_unikernel_0__dout),
    .t1_s_empty_n(k_rd_unikernel_0__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_0__empty_n),
    .t1_s_read(k_rd_unikernel_0__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_0__din),
    .t0_full_n(k_wr_unikernel_0__full_n),
    .t0_write(k_wr_unikernel_0__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_1__ap_start),
    .ap_done(JACOBI3D_1__ap_done),
    .ap_idle(JACOBI3D_1__ap_idle),
    .ap_ready(JACOBI3D_1__ap_ready),
    .iters(JACOBI3D_1___iters__q0),
    .t1_s_dout(k_rd_unikernel_1__dout),
    .t1_peek_dout(k_rd_unikernel_1__dout),
    .t1_s_empty_n(k_rd_unikernel_1__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_1__empty_n),
    .t1_s_read(k_rd_unikernel_1__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_1__din),
    .t0_full_n(k_wr_unikernel_1__full_n),
    .t0_write(k_wr_unikernel_1__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_2__ap_start),
    .ap_done(JACOBI3D_2__ap_done),
    .ap_idle(JACOBI3D_2__ap_idle),
    .ap_ready(JACOBI3D_2__ap_ready),
    .iters(JACOBI3D_2___iters__q0),
    .t1_s_dout(k_rd_unikernel_2__dout),
    .t1_peek_dout(k_rd_unikernel_2__dout),
    .t1_s_empty_n(k_rd_unikernel_2__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_2__empty_n),
    .t1_s_read(k_rd_unikernel_2__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_2__din),
    .t0_full_n(k_wr_unikernel_2__full_n),
    .t0_write(k_wr_unikernel_2__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_3__ap_start),
    .ap_done(JACOBI3D_3__ap_done),
    .ap_idle(JACOBI3D_3__ap_idle),
    .ap_ready(JACOBI3D_3__ap_ready),
    .iters(JACOBI3D_3___iters__q0),
    .t1_s_dout(k_rd_unikernel_3__dout),
    .t1_peek_dout(k_rd_unikernel_3__dout),
    .t1_s_empty_n(k_rd_unikernel_3__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_3__empty_n),
    .t1_s_read(k_rd_unikernel_3__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_3__din),
    .t0_full_n(k_wr_unikernel_3__full_n),
    .t0_write(k_wr_unikernel_3__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_4__ap_start),
    .ap_done(JACOBI3D_4__ap_done),
    .ap_idle(JACOBI3D_4__ap_idle),
    .ap_ready(JACOBI3D_4__ap_ready),
    .iters(JACOBI3D_4___iters__q0),
    .t1_s_dout(k_rd_unikernel_4__dout),
    .t1_peek_dout(k_rd_unikernel_4__dout),
    .t1_s_empty_n(k_rd_unikernel_4__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_4__empty_n),
    .t1_s_read(k_rd_unikernel_4__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_4__din),
    .t0_full_n(k_wr_unikernel_4__full_n),
    .t0_write(k_wr_unikernel_4__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_5__ap_start),
    .ap_done(JACOBI3D_5__ap_done),
    .ap_idle(JACOBI3D_5__ap_idle),
    .ap_ready(JACOBI3D_5__ap_ready),
    .iters(JACOBI3D_5___iters__q0),
    .t1_s_dout(k_rd_unikernel_5__dout),
    .t1_peek_dout(k_rd_unikernel_5__dout),
    .t1_s_empty_n(k_rd_unikernel_5__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_5__empty_n),
    .t1_s_read(k_rd_unikernel_5__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_5__din),
    .t0_full_n(k_wr_unikernel_5__full_n),
    .t0_write(k_wr_unikernel_5__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_6__ap_start),
    .ap_done(JACOBI3D_6__ap_done),
    .ap_idle(JACOBI3D_6__ap_idle),
    .ap_ready(JACOBI3D_6__ap_ready),
    .iters(JACOBI3D_6___iters__q0),
    .t1_s_dout(k_rd_unikernel_6__dout),
    .t1_peek_dout(k_rd_unikernel_6__dout),
    .t1_s_empty_n(k_rd_unikernel_6__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_6__empty_n),
    .t1_s_read(k_rd_unikernel_6__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_6__din),
    .t0_full_n(k_wr_unikernel_6__full_n),
    .t0_write(k_wr_unikernel_6__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_7__ap_start),
    .ap_done(JACOBI3D_7__ap_done),
    .ap_idle(JACOBI3D_7__ap_idle),
    .ap_ready(JACOBI3D_7__ap_ready),
    .iters(JACOBI3D_7___iters__q0),
    .t1_s_dout(k_rd_unikernel_7__dout),
    .t1_peek_dout(k_rd_unikernel_7__dout),
    .t1_s_empty_n(k_rd_unikernel_7__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_7__empty_n),
    .t1_s_read(k_rd_unikernel_7__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_7__din),
    .t0_full_n(k_wr_unikernel_7__full_n),
    .t0_write(k_wr_unikernel_7__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_8__ap_start),
    .ap_done(JACOBI3D_8__ap_done),
    .ap_idle(JACOBI3D_8__ap_idle),
    .ap_ready(JACOBI3D_8__ap_ready),
    .iters(JACOBI3D_8___iters__q0),
    .t1_s_dout(k_rd_unikernel_8__dout),
    .t1_peek_dout(k_rd_unikernel_8__dout),
    .t1_s_empty_n(k_rd_unikernel_8__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_8__empty_n),
    .t1_s_read(k_rd_unikernel_8__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_8__din),
    .t0_full_n(k_wr_unikernel_8__full_n),
    .t0_write(k_wr_unikernel_8__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_9__ap_start),
    .ap_done(JACOBI3D_9__ap_done),
    .ap_idle(JACOBI3D_9__ap_idle),
    .ap_ready(JACOBI3D_9__ap_ready),
    .iters(JACOBI3D_9___iters__q0),
    .t1_s_dout(k_rd_unikernel_9__dout),
    .t1_peek_dout(k_rd_unikernel_9__dout),
    .t1_s_empty_n(k_rd_unikernel_9__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_9__empty_n),
    .t1_s_read(k_rd_unikernel_9__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_9__din),
    .t0_full_n(k_wr_unikernel_9__full_n),
    .t0_write(k_wr_unikernel_9__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_10__ap_start),
    .ap_done(JACOBI3D_10__ap_done),
    .ap_idle(JACOBI3D_10__ap_idle),
    .ap_ready(JACOBI3D_10__ap_ready),
    .iters(JACOBI3D_10___iters__q0),
    .t1_s_dout(k_rd_unikernel_10__dout),
    .t1_peek_dout(k_rd_unikernel_10__dout),
    .t1_s_empty_n(k_rd_unikernel_10__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_10__empty_n),
    .t1_s_read(k_rd_unikernel_10__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_10__din),
    .t0_full_n(k_wr_unikernel_10__full_n),
    .t0_write(k_wr_unikernel_10__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_11__ap_start),
    .ap_done(JACOBI3D_11__ap_done),
    .ap_idle(JACOBI3D_11__ap_idle),
    .ap_ready(JACOBI3D_11__ap_ready),
    .iters(JACOBI3D_11___iters__q0),
    .t1_s_dout(k_rd_unikernel_11__dout),
    .t1_peek_dout(k_rd_unikernel_11__dout),
    .t1_s_empty_n(k_rd_unikernel_11__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_11__empty_n),
    .t1_s_read(k_rd_unikernel_11__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_11__din),
    .t0_full_n(k_wr_unikernel_11__full_n),
    .t0_write(k_wr_unikernel_11__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_12__ap_start),
    .ap_done(JACOBI3D_12__ap_done),
    .ap_idle(JACOBI3D_12__ap_idle),
    .ap_ready(JACOBI3D_12__ap_ready),
    .iters(JACOBI3D_12___iters__q0),
    .t1_s_dout(k_rd_unikernel_12__dout),
    .t1_peek_dout(k_rd_unikernel_12__dout),
    .t1_s_empty_n(k_rd_unikernel_12__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_12__empty_n),
    .t1_s_read(k_rd_unikernel_12__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_12__din),
    .t0_full_n(k_wr_unikernel_12__full_n),
    .t0_write(k_wr_unikernel_12__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_13__ap_start),
    .ap_done(JACOBI3D_13__ap_done),
    .ap_idle(JACOBI3D_13__ap_idle),
    .ap_ready(JACOBI3D_13__ap_ready),
    .iters(JACOBI3D_13___iters__q0),
    .t1_s_dout(k_rd_unikernel_13__dout),
    .t1_peek_dout(k_rd_unikernel_13__dout),
    .t1_s_empty_n(k_rd_unikernel_13__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_13__empty_n),
    .t1_s_read(k_rd_unikernel_13__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_13__din),
    .t0_full_n(k_wr_unikernel_13__full_n),
    .t0_write(k_wr_unikernel_13__write)
  );


  (* keep_hierarchy = "yes" *) JACOBI3D
  JACOBI3D_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(JACOBI3D_14__ap_start),
    .ap_done(JACOBI3D_14__ap_done),
    .ap_idle(JACOBI3D_14__ap_idle),
    .ap_ready(JACOBI3D_14__ap_ready),
    .iters(JACOBI3D_14___iters__q0),
    .t1_s_dout(k_rd_unikernel_14__dout),
    .t1_peek_dout(k_rd_unikernel_14__dout),
    .t1_s_empty_n(k_rd_unikernel_14__empty_n),
    .t1_peek_empty_n(k_rd_unikernel_14__empty_n),
    .t1_s_read(k_rd_unikernel_14__read),
    .t1_peek_read(),
    .t0_din(k_wr_unikernel_14__din),
    .t0_full_n(k_wr_unikernel_14__full_n),
    .t0_write(k_wr_unikernel_14__write)
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_0__ap_start),
    .ap_done(inter_kernel_0__ap_done),
    .ap_idle(inter_kernel_0__ap_idle),
    .ap_ready(inter_kernel_0__ap_ready),
    .a_read_addr_din(in_0_read_addr__din),
    .a_read_addr_full_n(in_0_read_addr__full_n),
    .a_read_addr_write(in_0_read_addr__write),
    .a_read_data_s_dout({1'b0, in_0_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_0_read_data__dout}),
    .a_read_data_s_empty_n(in_0_read_data__empty_n),
    .a_read_data_peek_empty_n(in_0_read_data__empty_n),
    .a_read_data_s_read(in_0_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_0_write_addr__din),
    .a_write_addr_full_n(in_0_write_addr__full_n),
    .a_write_addr_write(in_0_write_addr__write),
    .a_write_data_din(in_0_write_data__din),
    .a_write_data_full_n(in_0_write_data__full_n),
    .a_write_data_write(in_0_write_data__write),
    .a_write_resp_s_dout({1'b0, in_0_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_0_write_resp__dout}),
    .a_write_resp_s_empty_n(in_0_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_0_write_resp__empty_n),
    .a_write_resp_s_read(in_0_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_0___iters__q0),
    .stream_out_din(k_rd_unikernel_0__din),
    .stream_out_full_n(k_rd_unikernel_0__full_n),
    .stream_out_write(k_rd_unikernel_0__write),
    .stream_in_s_dout(k_wr_unikernel_0__dout),
    .stream_in_peek_dout(k_wr_unikernel_0__dout),
    .stream_in_s_empty_n(k_wr_unikernel_0__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_0__empty_n),
    .stream_in_s_read(k_wr_unikernel_0__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_0_read_addr__din),
    .b_read_addr_full_n(out_0_read_addr__full_n),
    .b_read_addr_write(out_0_read_addr__write),
    .b_read_data_s_dout({1'b0, out_0_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_0_read_data__dout}),
    .b_read_data_s_empty_n(out_0_read_data__empty_n),
    .b_read_data_peek_empty_n(out_0_read_data__empty_n),
    .b_read_data_s_read(out_0_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_0_write_addr__din),
    .b_write_addr_full_n(out_0_write_addr__full_n),
    .b_write_addr_write(out_0_write_addr__write),
    .b_write_data_din(out_0_write_data__din),
    .b_write_data_full_n(out_0_write_data__full_n),
    .b_write_data_write(out_0_write_data__write),
    .b_write_resp_s_dout({1'b0, out_0_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_0_write_resp__dout}),
    .b_write_resp_s_empty_n(out_0_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_0_write_resp__empty_n),
    .b_write_resp_s_read(out_0_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_1__ap_start),
    .ap_done(inter_kernel_1__ap_done),
    .ap_idle(inter_kernel_1__ap_idle),
    .ap_ready(inter_kernel_1__ap_ready),
    .a_read_addr_din(in_1_read_addr__din),
    .a_read_addr_full_n(in_1_read_addr__full_n),
    .a_read_addr_write(in_1_read_addr__write),
    .a_read_data_s_dout({1'b0, in_1_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_1_read_data__dout}),
    .a_read_data_s_empty_n(in_1_read_data__empty_n),
    .a_read_data_peek_empty_n(in_1_read_data__empty_n),
    .a_read_data_s_read(in_1_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_1_write_addr__din),
    .a_write_addr_full_n(in_1_write_addr__full_n),
    .a_write_addr_write(in_1_write_addr__write),
    .a_write_data_din(in_1_write_data__din),
    .a_write_data_full_n(in_1_write_data__full_n),
    .a_write_data_write(in_1_write_data__write),
    .a_write_resp_s_dout({1'b0, in_1_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_1_write_resp__dout}),
    .a_write_resp_s_empty_n(in_1_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_1_write_resp__empty_n),
    .a_write_resp_s_read(in_1_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_1___iters__q0),
    .stream_out_din(k_rd_unikernel_1__din),
    .stream_out_full_n(k_rd_unikernel_1__full_n),
    .stream_out_write(k_rd_unikernel_1__write),
    .stream_in_s_dout(k_wr_unikernel_1__dout),
    .stream_in_peek_dout(k_wr_unikernel_1__dout),
    .stream_in_s_empty_n(k_wr_unikernel_1__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_1__empty_n),
    .stream_in_s_read(k_wr_unikernel_1__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_1_read_addr__din),
    .b_read_addr_full_n(out_1_read_addr__full_n),
    .b_read_addr_write(out_1_read_addr__write),
    .b_read_data_s_dout({1'b0, out_1_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_1_read_data__dout}),
    .b_read_data_s_empty_n(out_1_read_data__empty_n),
    .b_read_data_peek_empty_n(out_1_read_data__empty_n),
    .b_read_data_s_read(out_1_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_1_write_addr__din),
    .b_write_addr_full_n(out_1_write_addr__full_n),
    .b_write_addr_write(out_1_write_addr__write),
    .b_write_data_din(out_1_write_data__din),
    .b_write_data_full_n(out_1_write_data__full_n),
    .b_write_data_write(out_1_write_data__write),
    .b_write_resp_s_dout({1'b0, out_1_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_1_write_resp__dout}),
    .b_write_resp_s_empty_n(out_1_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_1_write_resp__empty_n),
    .b_write_resp_s_read(out_1_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_2__ap_start),
    .ap_done(inter_kernel_2__ap_done),
    .ap_idle(inter_kernel_2__ap_idle),
    .ap_ready(inter_kernel_2__ap_ready),
    .a_read_addr_din(in_2_read_addr__din),
    .a_read_addr_full_n(in_2_read_addr__full_n),
    .a_read_addr_write(in_2_read_addr__write),
    .a_read_data_s_dout({1'b0, in_2_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_2_read_data__dout}),
    .a_read_data_s_empty_n(in_2_read_data__empty_n),
    .a_read_data_peek_empty_n(in_2_read_data__empty_n),
    .a_read_data_s_read(in_2_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_2_write_addr__din),
    .a_write_addr_full_n(in_2_write_addr__full_n),
    .a_write_addr_write(in_2_write_addr__write),
    .a_write_data_din(in_2_write_data__din),
    .a_write_data_full_n(in_2_write_data__full_n),
    .a_write_data_write(in_2_write_data__write),
    .a_write_resp_s_dout({1'b0, in_2_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_2_write_resp__dout}),
    .a_write_resp_s_empty_n(in_2_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_2_write_resp__empty_n),
    .a_write_resp_s_read(in_2_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_2___iters__q0),
    .stream_out_din(k_rd_unikernel_2__din),
    .stream_out_full_n(k_rd_unikernel_2__full_n),
    .stream_out_write(k_rd_unikernel_2__write),
    .stream_in_s_dout(k_wr_unikernel_2__dout),
    .stream_in_peek_dout(k_wr_unikernel_2__dout),
    .stream_in_s_empty_n(k_wr_unikernel_2__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_2__empty_n),
    .stream_in_s_read(k_wr_unikernel_2__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_2_read_addr__din),
    .b_read_addr_full_n(out_2_read_addr__full_n),
    .b_read_addr_write(out_2_read_addr__write),
    .b_read_data_s_dout({1'b0, out_2_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_2_read_data__dout}),
    .b_read_data_s_empty_n(out_2_read_data__empty_n),
    .b_read_data_peek_empty_n(out_2_read_data__empty_n),
    .b_read_data_s_read(out_2_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_2_write_addr__din),
    .b_write_addr_full_n(out_2_write_addr__full_n),
    .b_write_addr_write(out_2_write_addr__write),
    .b_write_data_din(out_2_write_data__din),
    .b_write_data_full_n(out_2_write_data__full_n),
    .b_write_data_write(out_2_write_data__write),
    .b_write_resp_s_dout({1'b0, out_2_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_2_write_resp__dout}),
    .b_write_resp_s_empty_n(out_2_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_2_write_resp__empty_n),
    .b_write_resp_s_read(out_2_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_3__ap_start),
    .ap_done(inter_kernel_3__ap_done),
    .ap_idle(inter_kernel_3__ap_idle),
    .ap_ready(inter_kernel_3__ap_ready),
    .a_read_addr_din(in_3_read_addr__din),
    .a_read_addr_full_n(in_3_read_addr__full_n),
    .a_read_addr_write(in_3_read_addr__write),
    .a_read_data_s_dout({1'b0, in_3_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_3_read_data__dout}),
    .a_read_data_s_empty_n(in_3_read_data__empty_n),
    .a_read_data_peek_empty_n(in_3_read_data__empty_n),
    .a_read_data_s_read(in_3_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_3_write_addr__din),
    .a_write_addr_full_n(in_3_write_addr__full_n),
    .a_write_addr_write(in_3_write_addr__write),
    .a_write_data_din(in_3_write_data__din),
    .a_write_data_full_n(in_3_write_data__full_n),
    .a_write_data_write(in_3_write_data__write),
    .a_write_resp_s_dout({1'b0, in_3_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_3_write_resp__dout}),
    .a_write_resp_s_empty_n(in_3_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_3_write_resp__empty_n),
    .a_write_resp_s_read(in_3_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_3___iters__q0),
    .stream_out_din(k_rd_unikernel_3__din),
    .stream_out_full_n(k_rd_unikernel_3__full_n),
    .stream_out_write(k_rd_unikernel_3__write),
    .stream_in_s_dout(k_wr_unikernel_3__dout),
    .stream_in_peek_dout(k_wr_unikernel_3__dout),
    .stream_in_s_empty_n(k_wr_unikernel_3__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_3__empty_n),
    .stream_in_s_read(k_wr_unikernel_3__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_3_read_addr__din),
    .b_read_addr_full_n(out_3_read_addr__full_n),
    .b_read_addr_write(out_3_read_addr__write),
    .b_read_data_s_dout({1'b0, out_3_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_3_read_data__dout}),
    .b_read_data_s_empty_n(out_3_read_data__empty_n),
    .b_read_data_peek_empty_n(out_3_read_data__empty_n),
    .b_read_data_s_read(out_3_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_3_write_addr__din),
    .b_write_addr_full_n(out_3_write_addr__full_n),
    .b_write_addr_write(out_3_write_addr__write),
    .b_write_data_din(out_3_write_data__din),
    .b_write_data_full_n(out_3_write_data__full_n),
    .b_write_data_write(out_3_write_data__write),
    .b_write_resp_s_dout({1'b0, out_3_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_3_write_resp__dout}),
    .b_write_resp_s_empty_n(out_3_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_3_write_resp__empty_n),
    .b_write_resp_s_read(out_3_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_4__ap_start),
    .ap_done(inter_kernel_4__ap_done),
    .ap_idle(inter_kernel_4__ap_idle),
    .ap_ready(inter_kernel_4__ap_ready),
    .a_read_addr_din(in_4_read_addr__din),
    .a_read_addr_full_n(in_4_read_addr__full_n),
    .a_read_addr_write(in_4_read_addr__write),
    .a_read_data_s_dout({1'b0, in_4_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_4_read_data__dout}),
    .a_read_data_s_empty_n(in_4_read_data__empty_n),
    .a_read_data_peek_empty_n(in_4_read_data__empty_n),
    .a_read_data_s_read(in_4_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_4_write_addr__din),
    .a_write_addr_full_n(in_4_write_addr__full_n),
    .a_write_addr_write(in_4_write_addr__write),
    .a_write_data_din(in_4_write_data__din),
    .a_write_data_full_n(in_4_write_data__full_n),
    .a_write_data_write(in_4_write_data__write),
    .a_write_resp_s_dout({1'b0, in_4_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_4_write_resp__dout}),
    .a_write_resp_s_empty_n(in_4_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_4_write_resp__empty_n),
    .a_write_resp_s_read(in_4_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_4___iters__q0),
    .stream_out_din(k_rd_unikernel_4__din),
    .stream_out_full_n(k_rd_unikernel_4__full_n),
    .stream_out_write(k_rd_unikernel_4__write),
    .stream_in_s_dout(k_wr_unikernel_4__dout),
    .stream_in_peek_dout(k_wr_unikernel_4__dout),
    .stream_in_s_empty_n(k_wr_unikernel_4__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_4__empty_n),
    .stream_in_s_read(k_wr_unikernel_4__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_4_read_addr__din),
    .b_read_addr_full_n(out_4_read_addr__full_n),
    .b_read_addr_write(out_4_read_addr__write),
    .b_read_data_s_dout({1'b0, out_4_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_4_read_data__dout}),
    .b_read_data_s_empty_n(out_4_read_data__empty_n),
    .b_read_data_peek_empty_n(out_4_read_data__empty_n),
    .b_read_data_s_read(out_4_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_4_write_addr__din),
    .b_write_addr_full_n(out_4_write_addr__full_n),
    .b_write_addr_write(out_4_write_addr__write),
    .b_write_data_din(out_4_write_data__din),
    .b_write_data_full_n(out_4_write_data__full_n),
    .b_write_data_write(out_4_write_data__write),
    .b_write_resp_s_dout({1'b0, out_4_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_4_write_resp__dout}),
    .b_write_resp_s_empty_n(out_4_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_4_write_resp__empty_n),
    .b_write_resp_s_read(out_4_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_5__ap_start),
    .ap_done(inter_kernel_5__ap_done),
    .ap_idle(inter_kernel_5__ap_idle),
    .ap_ready(inter_kernel_5__ap_ready),
    .a_read_addr_din(in_5_read_addr__din),
    .a_read_addr_full_n(in_5_read_addr__full_n),
    .a_read_addr_write(in_5_read_addr__write),
    .a_read_data_s_dout({1'b0, in_5_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_5_read_data__dout}),
    .a_read_data_s_empty_n(in_5_read_data__empty_n),
    .a_read_data_peek_empty_n(in_5_read_data__empty_n),
    .a_read_data_s_read(in_5_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_5_write_addr__din),
    .a_write_addr_full_n(in_5_write_addr__full_n),
    .a_write_addr_write(in_5_write_addr__write),
    .a_write_data_din(in_5_write_data__din),
    .a_write_data_full_n(in_5_write_data__full_n),
    .a_write_data_write(in_5_write_data__write),
    .a_write_resp_s_dout({1'b0, in_5_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_5_write_resp__dout}),
    .a_write_resp_s_empty_n(in_5_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_5_write_resp__empty_n),
    .a_write_resp_s_read(in_5_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_5___iters__q0),
    .stream_out_din(k_rd_unikernel_5__din),
    .stream_out_full_n(k_rd_unikernel_5__full_n),
    .stream_out_write(k_rd_unikernel_5__write),
    .stream_in_s_dout(k_wr_unikernel_5__dout),
    .stream_in_peek_dout(k_wr_unikernel_5__dout),
    .stream_in_s_empty_n(k_wr_unikernel_5__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_5__empty_n),
    .stream_in_s_read(k_wr_unikernel_5__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_5_read_addr__din),
    .b_read_addr_full_n(out_5_read_addr__full_n),
    .b_read_addr_write(out_5_read_addr__write),
    .b_read_data_s_dout({1'b0, out_5_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_5_read_data__dout}),
    .b_read_data_s_empty_n(out_5_read_data__empty_n),
    .b_read_data_peek_empty_n(out_5_read_data__empty_n),
    .b_read_data_s_read(out_5_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_5_write_addr__din),
    .b_write_addr_full_n(out_5_write_addr__full_n),
    .b_write_addr_write(out_5_write_addr__write),
    .b_write_data_din(out_5_write_data__din),
    .b_write_data_full_n(out_5_write_data__full_n),
    .b_write_data_write(out_5_write_data__write),
    .b_write_resp_s_dout({1'b0, out_5_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_5_write_resp__dout}),
    .b_write_resp_s_empty_n(out_5_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_5_write_resp__empty_n),
    .b_write_resp_s_read(out_5_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_6__ap_start),
    .ap_done(inter_kernel_6__ap_done),
    .ap_idle(inter_kernel_6__ap_idle),
    .ap_ready(inter_kernel_6__ap_ready),
    .a_read_addr_din(in_6_read_addr__din),
    .a_read_addr_full_n(in_6_read_addr__full_n),
    .a_read_addr_write(in_6_read_addr__write),
    .a_read_data_s_dout({1'b0, in_6_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_6_read_data__dout}),
    .a_read_data_s_empty_n(in_6_read_data__empty_n),
    .a_read_data_peek_empty_n(in_6_read_data__empty_n),
    .a_read_data_s_read(in_6_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_6_write_addr__din),
    .a_write_addr_full_n(in_6_write_addr__full_n),
    .a_write_addr_write(in_6_write_addr__write),
    .a_write_data_din(in_6_write_data__din),
    .a_write_data_full_n(in_6_write_data__full_n),
    .a_write_data_write(in_6_write_data__write),
    .a_write_resp_s_dout({1'b0, in_6_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_6_write_resp__dout}),
    .a_write_resp_s_empty_n(in_6_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_6_write_resp__empty_n),
    .a_write_resp_s_read(in_6_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_6___iters__q0),
    .stream_out_din(k_rd_unikernel_6__din),
    .stream_out_full_n(k_rd_unikernel_6__full_n),
    .stream_out_write(k_rd_unikernel_6__write),
    .stream_in_s_dout(k_wr_unikernel_6__dout),
    .stream_in_peek_dout(k_wr_unikernel_6__dout),
    .stream_in_s_empty_n(k_wr_unikernel_6__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_6__empty_n),
    .stream_in_s_read(k_wr_unikernel_6__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_6_read_addr__din),
    .b_read_addr_full_n(out_6_read_addr__full_n),
    .b_read_addr_write(out_6_read_addr__write),
    .b_read_data_s_dout({1'b0, out_6_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_6_read_data__dout}),
    .b_read_data_s_empty_n(out_6_read_data__empty_n),
    .b_read_data_peek_empty_n(out_6_read_data__empty_n),
    .b_read_data_s_read(out_6_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_6_write_addr__din),
    .b_write_addr_full_n(out_6_write_addr__full_n),
    .b_write_addr_write(out_6_write_addr__write),
    .b_write_data_din(out_6_write_data__din),
    .b_write_data_full_n(out_6_write_data__full_n),
    .b_write_data_write(out_6_write_data__write),
    .b_write_resp_s_dout({1'b0, out_6_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_6_write_resp__dout}),
    .b_write_resp_s_empty_n(out_6_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_6_write_resp__empty_n),
    .b_write_resp_s_read(out_6_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_7__ap_start),
    .ap_done(inter_kernel_7__ap_done),
    .ap_idle(inter_kernel_7__ap_idle),
    .ap_ready(inter_kernel_7__ap_ready),
    .a_read_addr_din(in_7_read_addr__din),
    .a_read_addr_full_n(in_7_read_addr__full_n),
    .a_read_addr_write(in_7_read_addr__write),
    .a_read_data_s_dout({1'b0, in_7_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_7_read_data__dout}),
    .a_read_data_s_empty_n(in_7_read_data__empty_n),
    .a_read_data_peek_empty_n(in_7_read_data__empty_n),
    .a_read_data_s_read(in_7_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_7_write_addr__din),
    .a_write_addr_full_n(in_7_write_addr__full_n),
    .a_write_addr_write(in_7_write_addr__write),
    .a_write_data_din(in_7_write_data__din),
    .a_write_data_full_n(in_7_write_data__full_n),
    .a_write_data_write(in_7_write_data__write),
    .a_write_resp_s_dout({1'b0, in_7_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_7_write_resp__dout}),
    .a_write_resp_s_empty_n(in_7_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_7_write_resp__empty_n),
    .a_write_resp_s_read(in_7_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_7___iters__q0),
    .stream_out_din(k_rd_unikernel_7__din),
    .stream_out_full_n(k_rd_unikernel_7__full_n),
    .stream_out_write(k_rd_unikernel_7__write),
    .stream_in_s_dout(k_wr_unikernel_7__dout),
    .stream_in_peek_dout(k_wr_unikernel_7__dout),
    .stream_in_s_empty_n(k_wr_unikernel_7__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_7__empty_n),
    .stream_in_s_read(k_wr_unikernel_7__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_7_read_addr__din),
    .b_read_addr_full_n(out_7_read_addr__full_n),
    .b_read_addr_write(out_7_read_addr__write),
    .b_read_data_s_dout({1'b0, out_7_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_7_read_data__dout}),
    .b_read_data_s_empty_n(out_7_read_data__empty_n),
    .b_read_data_peek_empty_n(out_7_read_data__empty_n),
    .b_read_data_s_read(out_7_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_7_write_addr__din),
    .b_write_addr_full_n(out_7_write_addr__full_n),
    .b_write_addr_write(out_7_write_addr__write),
    .b_write_data_din(out_7_write_data__din),
    .b_write_data_full_n(out_7_write_data__full_n),
    .b_write_data_write(out_7_write_data__write),
    .b_write_resp_s_dout({1'b0, out_7_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_7_write_resp__dout}),
    .b_write_resp_s_empty_n(out_7_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_7_write_resp__empty_n),
    .b_write_resp_s_read(out_7_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_8__ap_start),
    .ap_done(inter_kernel_8__ap_done),
    .ap_idle(inter_kernel_8__ap_idle),
    .ap_ready(inter_kernel_8__ap_ready),
    .a_read_addr_din(in_8_read_addr__din),
    .a_read_addr_full_n(in_8_read_addr__full_n),
    .a_read_addr_write(in_8_read_addr__write),
    .a_read_data_s_dout({1'b0, in_8_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_8_read_data__dout}),
    .a_read_data_s_empty_n(in_8_read_data__empty_n),
    .a_read_data_peek_empty_n(in_8_read_data__empty_n),
    .a_read_data_s_read(in_8_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_8_write_addr__din),
    .a_write_addr_full_n(in_8_write_addr__full_n),
    .a_write_addr_write(in_8_write_addr__write),
    .a_write_data_din(in_8_write_data__din),
    .a_write_data_full_n(in_8_write_data__full_n),
    .a_write_data_write(in_8_write_data__write),
    .a_write_resp_s_dout({1'b0, in_8_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_8_write_resp__dout}),
    .a_write_resp_s_empty_n(in_8_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_8_write_resp__empty_n),
    .a_write_resp_s_read(in_8_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_8___iters__q0),
    .stream_out_din(k_rd_unikernel_8__din),
    .stream_out_full_n(k_rd_unikernel_8__full_n),
    .stream_out_write(k_rd_unikernel_8__write),
    .stream_in_s_dout(k_wr_unikernel_8__dout),
    .stream_in_peek_dout(k_wr_unikernel_8__dout),
    .stream_in_s_empty_n(k_wr_unikernel_8__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_8__empty_n),
    .stream_in_s_read(k_wr_unikernel_8__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_8_read_addr__din),
    .b_read_addr_full_n(out_8_read_addr__full_n),
    .b_read_addr_write(out_8_read_addr__write),
    .b_read_data_s_dout({1'b0, out_8_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_8_read_data__dout}),
    .b_read_data_s_empty_n(out_8_read_data__empty_n),
    .b_read_data_peek_empty_n(out_8_read_data__empty_n),
    .b_read_data_s_read(out_8_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_8_write_addr__din),
    .b_write_addr_full_n(out_8_write_addr__full_n),
    .b_write_addr_write(out_8_write_addr__write),
    .b_write_data_din(out_8_write_data__din),
    .b_write_data_full_n(out_8_write_data__full_n),
    .b_write_data_write(out_8_write_data__write),
    .b_write_resp_s_dout({1'b0, out_8_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_8_write_resp__dout}),
    .b_write_resp_s_empty_n(out_8_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_8_write_resp__empty_n),
    .b_write_resp_s_read(out_8_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_9__ap_start),
    .ap_done(inter_kernel_9__ap_done),
    .ap_idle(inter_kernel_9__ap_idle),
    .ap_ready(inter_kernel_9__ap_ready),
    .a_read_addr_din(in_9_read_addr__din),
    .a_read_addr_full_n(in_9_read_addr__full_n),
    .a_read_addr_write(in_9_read_addr__write),
    .a_read_data_s_dout({1'b0, in_9_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_9_read_data__dout}),
    .a_read_data_s_empty_n(in_9_read_data__empty_n),
    .a_read_data_peek_empty_n(in_9_read_data__empty_n),
    .a_read_data_s_read(in_9_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_9_write_addr__din),
    .a_write_addr_full_n(in_9_write_addr__full_n),
    .a_write_addr_write(in_9_write_addr__write),
    .a_write_data_din(in_9_write_data__din),
    .a_write_data_full_n(in_9_write_data__full_n),
    .a_write_data_write(in_9_write_data__write),
    .a_write_resp_s_dout({1'b0, in_9_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_9_write_resp__dout}),
    .a_write_resp_s_empty_n(in_9_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_9_write_resp__empty_n),
    .a_write_resp_s_read(in_9_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_9___iters__q0),
    .stream_out_din(k_rd_unikernel_9__din),
    .stream_out_full_n(k_rd_unikernel_9__full_n),
    .stream_out_write(k_rd_unikernel_9__write),
    .stream_in_s_dout(k_wr_unikernel_9__dout),
    .stream_in_peek_dout(k_wr_unikernel_9__dout),
    .stream_in_s_empty_n(k_wr_unikernel_9__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_9__empty_n),
    .stream_in_s_read(k_wr_unikernel_9__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_9_read_addr__din),
    .b_read_addr_full_n(out_9_read_addr__full_n),
    .b_read_addr_write(out_9_read_addr__write),
    .b_read_data_s_dout({1'b0, out_9_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_9_read_data__dout}),
    .b_read_data_s_empty_n(out_9_read_data__empty_n),
    .b_read_data_peek_empty_n(out_9_read_data__empty_n),
    .b_read_data_s_read(out_9_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_9_write_addr__din),
    .b_write_addr_full_n(out_9_write_addr__full_n),
    .b_write_addr_write(out_9_write_addr__write),
    .b_write_data_din(out_9_write_data__din),
    .b_write_data_full_n(out_9_write_data__full_n),
    .b_write_data_write(out_9_write_data__write),
    .b_write_resp_s_dout({1'b0, out_9_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_9_write_resp__dout}),
    .b_write_resp_s_empty_n(out_9_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_9_write_resp__empty_n),
    .b_write_resp_s_read(out_9_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_10__ap_start),
    .ap_done(inter_kernel_10__ap_done),
    .ap_idle(inter_kernel_10__ap_idle),
    .ap_ready(inter_kernel_10__ap_ready),
    .a_read_addr_din(in_10_read_addr__din),
    .a_read_addr_full_n(in_10_read_addr__full_n),
    .a_read_addr_write(in_10_read_addr__write),
    .a_read_data_s_dout({1'b0, in_10_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_10_read_data__dout}),
    .a_read_data_s_empty_n(in_10_read_data__empty_n),
    .a_read_data_peek_empty_n(in_10_read_data__empty_n),
    .a_read_data_s_read(in_10_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_10_write_addr__din),
    .a_write_addr_full_n(in_10_write_addr__full_n),
    .a_write_addr_write(in_10_write_addr__write),
    .a_write_data_din(in_10_write_data__din),
    .a_write_data_full_n(in_10_write_data__full_n),
    .a_write_data_write(in_10_write_data__write),
    .a_write_resp_s_dout({1'b0, in_10_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_10_write_resp__dout}),
    .a_write_resp_s_empty_n(in_10_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_10_write_resp__empty_n),
    .a_write_resp_s_read(in_10_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_10___iters__q0),
    .stream_out_din(k_rd_unikernel_10__din),
    .stream_out_full_n(k_rd_unikernel_10__full_n),
    .stream_out_write(k_rd_unikernel_10__write),
    .stream_in_s_dout(k_wr_unikernel_10__dout),
    .stream_in_peek_dout(k_wr_unikernel_10__dout),
    .stream_in_s_empty_n(k_wr_unikernel_10__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_10__empty_n),
    .stream_in_s_read(k_wr_unikernel_10__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_10_read_addr__din),
    .b_read_addr_full_n(out_10_read_addr__full_n),
    .b_read_addr_write(out_10_read_addr__write),
    .b_read_data_s_dout({1'b0, out_10_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_10_read_data__dout}),
    .b_read_data_s_empty_n(out_10_read_data__empty_n),
    .b_read_data_peek_empty_n(out_10_read_data__empty_n),
    .b_read_data_s_read(out_10_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_10_write_addr__din),
    .b_write_addr_full_n(out_10_write_addr__full_n),
    .b_write_addr_write(out_10_write_addr__write),
    .b_write_data_din(out_10_write_data__din),
    .b_write_data_full_n(out_10_write_data__full_n),
    .b_write_data_write(out_10_write_data__write),
    .b_write_resp_s_dout({1'b0, out_10_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_10_write_resp__dout}),
    .b_write_resp_s_empty_n(out_10_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_10_write_resp__empty_n),
    .b_write_resp_s_read(out_10_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_11__ap_start),
    .ap_done(inter_kernel_11__ap_done),
    .ap_idle(inter_kernel_11__ap_idle),
    .ap_ready(inter_kernel_11__ap_ready),
    .a_read_addr_din(in_11_read_addr__din),
    .a_read_addr_full_n(in_11_read_addr__full_n),
    .a_read_addr_write(in_11_read_addr__write),
    .a_read_data_s_dout({1'b0, in_11_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_11_read_data__dout}),
    .a_read_data_s_empty_n(in_11_read_data__empty_n),
    .a_read_data_peek_empty_n(in_11_read_data__empty_n),
    .a_read_data_s_read(in_11_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_11_write_addr__din),
    .a_write_addr_full_n(in_11_write_addr__full_n),
    .a_write_addr_write(in_11_write_addr__write),
    .a_write_data_din(in_11_write_data__din),
    .a_write_data_full_n(in_11_write_data__full_n),
    .a_write_data_write(in_11_write_data__write),
    .a_write_resp_s_dout({1'b0, in_11_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_11_write_resp__dout}),
    .a_write_resp_s_empty_n(in_11_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_11_write_resp__empty_n),
    .a_write_resp_s_read(in_11_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_11___iters__q0),
    .stream_out_din(k_rd_unikernel_11__din),
    .stream_out_full_n(k_rd_unikernel_11__full_n),
    .stream_out_write(k_rd_unikernel_11__write),
    .stream_in_s_dout(k_wr_unikernel_11__dout),
    .stream_in_peek_dout(k_wr_unikernel_11__dout),
    .stream_in_s_empty_n(k_wr_unikernel_11__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_11__empty_n),
    .stream_in_s_read(k_wr_unikernel_11__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_11_read_addr__din),
    .b_read_addr_full_n(out_11_read_addr__full_n),
    .b_read_addr_write(out_11_read_addr__write),
    .b_read_data_s_dout({1'b0, out_11_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_11_read_data__dout}),
    .b_read_data_s_empty_n(out_11_read_data__empty_n),
    .b_read_data_peek_empty_n(out_11_read_data__empty_n),
    .b_read_data_s_read(out_11_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_11_write_addr__din),
    .b_write_addr_full_n(out_11_write_addr__full_n),
    .b_write_addr_write(out_11_write_addr__write),
    .b_write_data_din(out_11_write_data__din),
    .b_write_data_full_n(out_11_write_data__full_n),
    .b_write_data_write(out_11_write_data__write),
    .b_write_resp_s_dout({1'b0, out_11_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_11_write_resp__dout}),
    .b_write_resp_s_empty_n(out_11_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_11_write_resp__empty_n),
    .b_write_resp_s_read(out_11_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_12__ap_start),
    .ap_done(inter_kernel_12__ap_done),
    .ap_idle(inter_kernel_12__ap_idle),
    .ap_ready(inter_kernel_12__ap_ready),
    .a_read_addr_din(in_12_read_addr__din),
    .a_read_addr_full_n(in_12_read_addr__full_n),
    .a_read_addr_write(in_12_read_addr__write),
    .a_read_data_s_dout({1'b0, in_12_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_12_read_data__dout}),
    .a_read_data_s_empty_n(in_12_read_data__empty_n),
    .a_read_data_peek_empty_n(in_12_read_data__empty_n),
    .a_read_data_s_read(in_12_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_12_write_addr__din),
    .a_write_addr_full_n(in_12_write_addr__full_n),
    .a_write_addr_write(in_12_write_addr__write),
    .a_write_data_din(in_12_write_data__din),
    .a_write_data_full_n(in_12_write_data__full_n),
    .a_write_data_write(in_12_write_data__write),
    .a_write_resp_s_dout({1'b0, in_12_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_12_write_resp__dout}),
    .a_write_resp_s_empty_n(in_12_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_12_write_resp__empty_n),
    .a_write_resp_s_read(in_12_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_12___iters__q0),
    .stream_out_din(k_rd_unikernel_12__din),
    .stream_out_full_n(k_rd_unikernel_12__full_n),
    .stream_out_write(k_rd_unikernel_12__write),
    .stream_in_s_dout(k_wr_unikernel_12__dout),
    .stream_in_peek_dout(k_wr_unikernel_12__dout),
    .stream_in_s_empty_n(k_wr_unikernel_12__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_12__empty_n),
    .stream_in_s_read(k_wr_unikernel_12__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_12_read_addr__din),
    .b_read_addr_full_n(out_12_read_addr__full_n),
    .b_read_addr_write(out_12_read_addr__write),
    .b_read_data_s_dout({1'b0, out_12_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_12_read_data__dout}),
    .b_read_data_s_empty_n(out_12_read_data__empty_n),
    .b_read_data_peek_empty_n(out_12_read_data__empty_n),
    .b_read_data_s_read(out_12_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_12_write_addr__din),
    .b_write_addr_full_n(out_12_write_addr__full_n),
    .b_write_addr_write(out_12_write_addr__write),
    .b_write_data_din(out_12_write_data__din),
    .b_write_data_full_n(out_12_write_data__full_n),
    .b_write_data_write(out_12_write_data__write),
    .b_write_resp_s_dout({1'b0, out_12_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_12_write_resp__dout}),
    .b_write_resp_s_empty_n(out_12_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_12_write_resp__empty_n),
    .b_write_resp_s_read(out_12_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_13__ap_start),
    .ap_done(inter_kernel_13__ap_done),
    .ap_idle(inter_kernel_13__ap_idle),
    .ap_ready(inter_kernel_13__ap_ready),
    .a_read_addr_din(in_13_read_addr__din),
    .a_read_addr_full_n(in_13_read_addr__full_n),
    .a_read_addr_write(in_13_read_addr__write),
    .a_read_data_s_dout({1'b0, in_13_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_13_read_data__dout}),
    .a_read_data_s_empty_n(in_13_read_data__empty_n),
    .a_read_data_peek_empty_n(in_13_read_data__empty_n),
    .a_read_data_s_read(in_13_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_13_write_addr__din),
    .a_write_addr_full_n(in_13_write_addr__full_n),
    .a_write_addr_write(in_13_write_addr__write),
    .a_write_data_din(in_13_write_data__din),
    .a_write_data_full_n(in_13_write_data__full_n),
    .a_write_data_write(in_13_write_data__write),
    .a_write_resp_s_dout({1'b0, in_13_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_13_write_resp__dout}),
    .a_write_resp_s_empty_n(in_13_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_13_write_resp__empty_n),
    .a_write_resp_s_read(in_13_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_13___iters__q0),
    .stream_out_din(k_rd_unikernel_13__din),
    .stream_out_full_n(k_rd_unikernel_13__full_n),
    .stream_out_write(k_rd_unikernel_13__write),
    .stream_in_s_dout(k_wr_unikernel_13__dout),
    .stream_in_peek_dout(k_wr_unikernel_13__dout),
    .stream_in_s_empty_n(k_wr_unikernel_13__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_13__empty_n),
    .stream_in_s_read(k_wr_unikernel_13__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_13_read_addr__din),
    .b_read_addr_full_n(out_13_read_addr__full_n),
    .b_read_addr_write(out_13_read_addr__write),
    .b_read_data_s_dout({1'b0, out_13_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_13_read_data__dout}),
    .b_read_data_s_empty_n(out_13_read_data__empty_n),
    .b_read_data_peek_empty_n(out_13_read_data__empty_n),
    .b_read_data_s_read(out_13_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_13_write_addr__din),
    .b_write_addr_full_n(out_13_write_addr__full_n),
    .b_write_addr_write(out_13_write_addr__write),
    .b_write_data_din(out_13_write_data__din),
    .b_write_data_full_n(out_13_write_data__full_n),
    .b_write_data_write(out_13_write_data__write),
    .b_write_resp_s_dout({1'b0, out_13_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_13_write_resp__dout}),
    .b_write_resp_s_empty_n(out_13_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_13_write_resp__empty_n),
    .b_write_resp_s_read(out_13_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) inter_kernel
  inter_kernel_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(inter_kernel_14__ap_start),
    .ap_done(inter_kernel_14__ap_done),
    .ap_idle(inter_kernel_14__ap_idle),
    .ap_ready(inter_kernel_14__ap_ready),
    .a_read_addr_din(in_14_read_addr__din),
    .a_read_addr_full_n(in_14_read_addr__full_n),
    .a_read_addr_write(in_14_read_addr__write),
    .a_read_data_s_dout({1'b0, in_14_read_data__dout}),
    .a_read_data_peek_dout({1'b0, in_14_read_data__dout}),
    .a_read_data_s_empty_n(in_14_read_data__empty_n),
    .a_read_data_peek_empty_n(in_14_read_data__empty_n),
    .a_read_data_s_read(in_14_read_data__read),
    .a_read_data_peek_read(),
    .a_write_addr_din(in_14_write_addr__din),
    .a_write_addr_full_n(in_14_write_addr__full_n),
    .a_write_addr_write(in_14_write_addr__write),
    .a_write_data_din(in_14_write_data__din),
    .a_write_data_full_n(in_14_write_data__full_n),
    .a_write_data_write(in_14_write_data__write),
    .a_write_resp_s_dout({1'b0, in_14_write_resp__dout}),
    .a_write_resp_peek_dout({1'b0, in_14_write_resp__dout}),
    .a_write_resp_s_empty_n(in_14_write_resp__empty_n),
    .a_write_resp_peek_empty_n(in_14_write_resp__empty_n),
    .a_write_resp_s_read(in_14_write_resp__read),
    .a_write_resp_peek_read(),
    .iters(inter_kernel_14___iters__q0),
    .stream_out_din(k_rd_unikernel_14__din),
    .stream_out_full_n(k_rd_unikernel_14__full_n),
    .stream_out_write(k_rd_unikernel_14__write),
    .stream_in_s_dout(k_wr_unikernel_14__dout),
    .stream_in_peek_dout(k_wr_unikernel_14__dout),
    .stream_in_s_empty_n(k_wr_unikernel_14__empty_n),
    .stream_in_peek_empty_n(k_wr_unikernel_14__empty_n),
    .stream_in_s_read(k_wr_unikernel_14__read),
    .stream_in_peek_read(),
    .b_read_addr_din(out_14_read_addr__din),
    .b_read_addr_full_n(out_14_read_addr__full_n),
    .b_read_addr_write(out_14_read_addr__write),
    .b_read_data_s_dout({1'b0, out_14_read_data__dout}),
    .b_read_data_peek_dout({1'b0, out_14_read_data__dout}),
    .b_read_data_s_empty_n(out_14_read_data__empty_n),
    .b_read_data_peek_empty_n(out_14_read_data__empty_n),
    .b_read_data_s_read(out_14_read_data__read),
    .b_read_data_peek_read(),
    .b_write_addr_din(out_14_write_addr__din),
    .b_write_addr_full_n(out_14_write_addr__full_n),
    .b_write_addr_write(out_14_write_addr__write),
    .b_write_data_din(out_14_write_data__din),
    .b_write_data_full_n(out_14_write_data__full_n),
    .b_write_data_write(out_14_write_data__write),
    .b_write_resp_s_dout({1'b0, out_14_write_resp__dout}),
    .b_write_resp_peek_dout({1'b0, out_14_write_resp__dout}),
    .b_write_resp_s_empty_n(out_14_write_resp__empty_n),
    .b_write_resp_peek_empty_n(out_14_write_resp__empty_n),
    .b_write_resp_s_read(out_14_write_resp__read),
    .b_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_0___in_0__q0),
    .m_axi_ARADDR(m_axi_in_0_ARADDR),
    .m_axi_ARBURST(m_axi_in_0_ARBURST),
    .m_axi_ARCACHE(m_axi_in_0_ARCACHE),
    .m_axi_ARID(m_axi_in_0_ARID),
    .m_axi_ARLEN(m_axi_in_0_ARLEN),
    .m_axi_ARLOCK(m_axi_in_0_ARLOCK),
    .m_axi_ARPROT(m_axi_in_0_ARPROT),
    .m_axi_ARQOS(m_axi_in_0_ARQOS),
    .m_axi_ARREADY(m_axi_in_0_ARREADY),
    .m_axi_ARSIZE(m_axi_in_0_ARSIZE),
    .m_axi_ARVALID(m_axi_in_0_ARVALID),
    .m_axi_AWADDR(m_axi_in_0_AWADDR),
    .m_axi_AWBURST(m_axi_in_0_AWBURST),
    .m_axi_AWCACHE(m_axi_in_0_AWCACHE),
    .m_axi_AWID(m_axi_in_0_AWID),
    .m_axi_AWLEN(m_axi_in_0_AWLEN),
    .m_axi_AWLOCK(m_axi_in_0_AWLOCK),
    .m_axi_AWPROT(m_axi_in_0_AWPROT),
    .m_axi_AWQOS(m_axi_in_0_AWQOS),
    .m_axi_AWREADY(m_axi_in_0_AWREADY),
    .m_axi_AWSIZE(m_axi_in_0_AWSIZE),
    .m_axi_AWVALID(m_axi_in_0_AWVALID),
    .m_axi_BID(m_axi_in_0_BID),
    .m_axi_BREADY(m_axi_in_0_BREADY),
    .m_axi_BRESP(m_axi_in_0_BRESP),
    .m_axi_BVALID(m_axi_in_0_BVALID),
    .m_axi_RDATA(m_axi_in_0_RDATA),
    .m_axi_RID(m_axi_in_0_RID),
    .m_axi_RLAST(m_axi_in_0_RLAST),
    .m_axi_RREADY(m_axi_in_0_RREADY),
    .m_axi_RRESP(m_axi_in_0_RRESP),
    .m_axi_RVALID(m_axi_in_0_RVALID),
    .m_axi_WDATA(m_axi_in_0_WDATA),
    .m_axi_WLAST(m_axi_in_0_WLAST),
    .m_axi_WREADY(m_axi_in_0_WREADY),
    .m_axi_WSTRB(m_axi_in_0_WSTRB),
    .m_axi_WVALID(m_axi_in_0_WVALID),
    .read_addr_din(in_0_read_addr__din),
    .read_addr_full_n(in_0_read_addr__full_n),
    .read_addr_write(in_0_read_addr__write),
    .read_data_dout(in_0_read_data__dout),
    .read_data_empty_n(in_0_read_data__empty_n),
    .read_data_read(in_0_read_data__read),
    .write_addr_din(in_0_write_addr__din),
    .write_addr_full_n(in_0_write_addr__full_n),
    .write_addr_write(in_0_write_addr__write),
    .write_data_din(in_0_write_data__din),
    .write_data_full_n(in_0_write_data__full_n),
    .write_data_write(in_0_write_data__write),
    .write_resp_dout(in_0_write_resp__dout),
    .write_resp_empty_n(in_0_write_resp__empty_n),
    .write_resp_read(in_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_0___out_0__q0),
    .m_axi_ARADDR(m_axi_out_0_ARADDR),
    .m_axi_ARBURST(m_axi_out_0_ARBURST),
    .m_axi_ARCACHE(m_axi_out_0_ARCACHE),
    .m_axi_ARID(m_axi_out_0_ARID),
    .m_axi_ARLEN(m_axi_out_0_ARLEN),
    .m_axi_ARLOCK(m_axi_out_0_ARLOCK),
    .m_axi_ARPROT(m_axi_out_0_ARPROT),
    .m_axi_ARQOS(m_axi_out_0_ARQOS),
    .m_axi_ARREADY(m_axi_out_0_ARREADY),
    .m_axi_ARSIZE(m_axi_out_0_ARSIZE),
    .m_axi_ARVALID(m_axi_out_0_ARVALID),
    .m_axi_AWADDR(m_axi_out_0_AWADDR),
    .m_axi_AWBURST(m_axi_out_0_AWBURST),
    .m_axi_AWCACHE(m_axi_out_0_AWCACHE),
    .m_axi_AWID(m_axi_out_0_AWID),
    .m_axi_AWLEN(m_axi_out_0_AWLEN),
    .m_axi_AWLOCK(m_axi_out_0_AWLOCK),
    .m_axi_AWPROT(m_axi_out_0_AWPROT),
    .m_axi_AWQOS(m_axi_out_0_AWQOS),
    .m_axi_AWREADY(m_axi_out_0_AWREADY),
    .m_axi_AWSIZE(m_axi_out_0_AWSIZE),
    .m_axi_AWVALID(m_axi_out_0_AWVALID),
    .m_axi_BID(m_axi_out_0_BID),
    .m_axi_BREADY(m_axi_out_0_BREADY),
    .m_axi_BRESP(m_axi_out_0_BRESP),
    .m_axi_BVALID(m_axi_out_0_BVALID),
    .m_axi_RDATA(m_axi_out_0_RDATA),
    .m_axi_RID(m_axi_out_0_RID),
    .m_axi_RLAST(m_axi_out_0_RLAST),
    .m_axi_RREADY(m_axi_out_0_RREADY),
    .m_axi_RRESP(m_axi_out_0_RRESP),
    .m_axi_RVALID(m_axi_out_0_RVALID),
    .m_axi_WDATA(m_axi_out_0_WDATA),
    .m_axi_WLAST(m_axi_out_0_WLAST),
    .m_axi_WREADY(m_axi_out_0_WREADY),
    .m_axi_WSTRB(m_axi_out_0_WSTRB),
    .m_axi_WVALID(m_axi_out_0_WVALID),
    .read_addr_din(out_0_read_addr__din),
    .read_addr_full_n(out_0_read_addr__full_n),
    .read_addr_write(out_0_read_addr__write),
    .read_data_dout(out_0_read_data__dout),
    .read_data_empty_n(out_0_read_data__empty_n),
    .read_data_read(out_0_read_data__read),
    .write_addr_din(out_0_write_addr__din),
    .write_addr_full_n(out_0_write_addr__full_n),
    .write_addr_write(out_0_write_addr__write),
    .write_data_din(out_0_write_data__din),
    .write_data_full_n(out_0_write_data__full_n),
    .write_data_write(out_0_write_data__write),
    .write_resp_dout(out_0_write_resp__dout),
    .write_resp_empty_n(out_0_write_resp__empty_n),
    .write_resp_read(out_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_1___in_1__q0),
    .m_axi_ARADDR(m_axi_in_1_ARADDR),
    .m_axi_ARBURST(m_axi_in_1_ARBURST),
    .m_axi_ARCACHE(m_axi_in_1_ARCACHE),
    .m_axi_ARID(m_axi_in_1_ARID),
    .m_axi_ARLEN(m_axi_in_1_ARLEN),
    .m_axi_ARLOCK(m_axi_in_1_ARLOCK),
    .m_axi_ARPROT(m_axi_in_1_ARPROT),
    .m_axi_ARQOS(m_axi_in_1_ARQOS),
    .m_axi_ARREADY(m_axi_in_1_ARREADY),
    .m_axi_ARSIZE(m_axi_in_1_ARSIZE),
    .m_axi_ARVALID(m_axi_in_1_ARVALID),
    .m_axi_AWADDR(m_axi_in_1_AWADDR),
    .m_axi_AWBURST(m_axi_in_1_AWBURST),
    .m_axi_AWCACHE(m_axi_in_1_AWCACHE),
    .m_axi_AWID(m_axi_in_1_AWID),
    .m_axi_AWLEN(m_axi_in_1_AWLEN),
    .m_axi_AWLOCK(m_axi_in_1_AWLOCK),
    .m_axi_AWPROT(m_axi_in_1_AWPROT),
    .m_axi_AWQOS(m_axi_in_1_AWQOS),
    .m_axi_AWREADY(m_axi_in_1_AWREADY),
    .m_axi_AWSIZE(m_axi_in_1_AWSIZE),
    .m_axi_AWVALID(m_axi_in_1_AWVALID),
    .m_axi_BID(m_axi_in_1_BID),
    .m_axi_BREADY(m_axi_in_1_BREADY),
    .m_axi_BRESP(m_axi_in_1_BRESP),
    .m_axi_BVALID(m_axi_in_1_BVALID),
    .m_axi_RDATA(m_axi_in_1_RDATA),
    .m_axi_RID(m_axi_in_1_RID),
    .m_axi_RLAST(m_axi_in_1_RLAST),
    .m_axi_RREADY(m_axi_in_1_RREADY),
    .m_axi_RRESP(m_axi_in_1_RRESP),
    .m_axi_RVALID(m_axi_in_1_RVALID),
    .m_axi_WDATA(m_axi_in_1_WDATA),
    .m_axi_WLAST(m_axi_in_1_WLAST),
    .m_axi_WREADY(m_axi_in_1_WREADY),
    .m_axi_WSTRB(m_axi_in_1_WSTRB),
    .m_axi_WVALID(m_axi_in_1_WVALID),
    .read_addr_din(in_1_read_addr__din),
    .read_addr_full_n(in_1_read_addr__full_n),
    .read_addr_write(in_1_read_addr__write),
    .read_data_dout(in_1_read_data__dout),
    .read_data_empty_n(in_1_read_data__empty_n),
    .read_data_read(in_1_read_data__read),
    .write_addr_din(in_1_write_addr__din),
    .write_addr_full_n(in_1_write_addr__full_n),
    .write_addr_write(in_1_write_addr__write),
    .write_data_din(in_1_write_data__din),
    .write_data_full_n(in_1_write_data__full_n),
    .write_data_write(in_1_write_data__write),
    .write_resp_dout(in_1_write_resp__dout),
    .write_resp_empty_n(in_1_write_resp__empty_n),
    .write_resp_read(in_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_1___out_1__q0),
    .m_axi_ARADDR(m_axi_out_1_ARADDR),
    .m_axi_ARBURST(m_axi_out_1_ARBURST),
    .m_axi_ARCACHE(m_axi_out_1_ARCACHE),
    .m_axi_ARID(m_axi_out_1_ARID),
    .m_axi_ARLEN(m_axi_out_1_ARLEN),
    .m_axi_ARLOCK(m_axi_out_1_ARLOCK),
    .m_axi_ARPROT(m_axi_out_1_ARPROT),
    .m_axi_ARQOS(m_axi_out_1_ARQOS),
    .m_axi_ARREADY(m_axi_out_1_ARREADY),
    .m_axi_ARSIZE(m_axi_out_1_ARSIZE),
    .m_axi_ARVALID(m_axi_out_1_ARVALID),
    .m_axi_AWADDR(m_axi_out_1_AWADDR),
    .m_axi_AWBURST(m_axi_out_1_AWBURST),
    .m_axi_AWCACHE(m_axi_out_1_AWCACHE),
    .m_axi_AWID(m_axi_out_1_AWID),
    .m_axi_AWLEN(m_axi_out_1_AWLEN),
    .m_axi_AWLOCK(m_axi_out_1_AWLOCK),
    .m_axi_AWPROT(m_axi_out_1_AWPROT),
    .m_axi_AWQOS(m_axi_out_1_AWQOS),
    .m_axi_AWREADY(m_axi_out_1_AWREADY),
    .m_axi_AWSIZE(m_axi_out_1_AWSIZE),
    .m_axi_AWVALID(m_axi_out_1_AWVALID),
    .m_axi_BID(m_axi_out_1_BID),
    .m_axi_BREADY(m_axi_out_1_BREADY),
    .m_axi_BRESP(m_axi_out_1_BRESP),
    .m_axi_BVALID(m_axi_out_1_BVALID),
    .m_axi_RDATA(m_axi_out_1_RDATA),
    .m_axi_RID(m_axi_out_1_RID),
    .m_axi_RLAST(m_axi_out_1_RLAST),
    .m_axi_RREADY(m_axi_out_1_RREADY),
    .m_axi_RRESP(m_axi_out_1_RRESP),
    .m_axi_RVALID(m_axi_out_1_RVALID),
    .m_axi_WDATA(m_axi_out_1_WDATA),
    .m_axi_WLAST(m_axi_out_1_WLAST),
    .m_axi_WREADY(m_axi_out_1_WREADY),
    .m_axi_WSTRB(m_axi_out_1_WSTRB),
    .m_axi_WVALID(m_axi_out_1_WVALID),
    .read_addr_din(out_1_read_addr__din),
    .read_addr_full_n(out_1_read_addr__full_n),
    .read_addr_write(out_1_read_addr__write),
    .read_data_dout(out_1_read_data__dout),
    .read_data_empty_n(out_1_read_data__empty_n),
    .read_data_read(out_1_read_data__read),
    .write_addr_din(out_1_write_addr__din),
    .write_addr_full_n(out_1_write_addr__full_n),
    .write_addr_write(out_1_write_addr__write),
    .write_data_din(out_1_write_data__din),
    .write_data_full_n(out_1_write_data__full_n),
    .write_data_write(out_1_write_data__write),
    .write_resp_dout(out_1_write_resp__dout),
    .write_resp_empty_n(out_1_write_resp__empty_n),
    .write_resp_read(out_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_2___in_2__q0),
    .m_axi_ARADDR(m_axi_in_2_ARADDR),
    .m_axi_ARBURST(m_axi_in_2_ARBURST),
    .m_axi_ARCACHE(m_axi_in_2_ARCACHE),
    .m_axi_ARID(m_axi_in_2_ARID),
    .m_axi_ARLEN(m_axi_in_2_ARLEN),
    .m_axi_ARLOCK(m_axi_in_2_ARLOCK),
    .m_axi_ARPROT(m_axi_in_2_ARPROT),
    .m_axi_ARQOS(m_axi_in_2_ARQOS),
    .m_axi_ARREADY(m_axi_in_2_ARREADY),
    .m_axi_ARSIZE(m_axi_in_2_ARSIZE),
    .m_axi_ARVALID(m_axi_in_2_ARVALID),
    .m_axi_AWADDR(m_axi_in_2_AWADDR),
    .m_axi_AWBURST(m_axi_in_2_AWBURST),
    .m_axi_AWCACHE(m_axi_in_2_AWCACHE),
    .m_axi_AWID(m_axi_in_2_AWID),
    .m_axi_AWLEN(m_axi_in_2_AWLEN),
    .m_axi_AWLOCK(m_axi_in_2_AWLOCK),
    .m_axi_AWPROT(m_axi_in_2_AWPROT),
    .m_axi_AWQOS(m_axi_in_2_AWQOS),
    .m_axi_AWREADY(m_axi_in_2_AWREADY),
    .m_axi_AWSIZE(m_axi_in_2_AWSIZE),
    .m_axi_AWVALID(m_axi_in_2_AWVALID),
    .m_axi_BID(m_axi_in_2_BID),
    .m_axi_BREADY(m_axi_in_2_BREADY),
    .m_axi_BRESP(m_axi_in_2_BRESP),
    .m_axi_BVALID(m_axi_in_2_BVALID),
    .m_axi_RDATA(m_axi_in_2_RDATA),
    .m_axi_RID(m_axi_in_2_RID),
    .m_axi_RLAST(m_axi_in_2_RLAST),
    .m_axi_RREADY(m_axi_in_2_RREADY),
    .m_axi_RRESP(m_axi_in_2_RRESP),
    .m_axi_RVALID(m_axi_in_2_RVALID),
    .m_axi_WDATA(m_axi_in_2_WDATA),
    .m_axi_WLAST(m_axi_in_2_WLAST),
    .m_axi_WREADY(m_axi_in_2_WREADY),
    .m_axi_WSTRB(m_axi_in_2_WSTRB),
    .m_axi_WVALID(m_axi_in_2_WVALID),
    .read_addr_din(in_2_read_addr__din),
    .read_addr_full_n(in_2_read_addr__full_n),
    .read_addr_write(in_2_read_addr__write),
    .read_data_dout(in_2_read_data__dout),
    .read_data_empty_n(in_2_read_data__empty_n),
    .read_data_read(in_2_read_data__read),
    .write_addr_din(in_2_write_addr__din),
    .write_addr_full_n(in_2_write_addr__full_n),
    .write_addr_write(in_2_write_addr__write),
    .write_data_din(in_2_write_data__din),
    .write_data_full_n(in_2_write_data__full_n),
    .write_data_write(in_2_write_data__write),
    .write_resp_dout(in_2_write_resp__dout),
    .write_resp_empty_n(in_2_write_resp__empty_n),
    .write_resp_read(in_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_2___out_2__q0),
    .m_axi_ARADDR(m_axi_out_2_ARADDR),
    .m_axi_ARBURST(m_axi_out_2_ARBURST),
    .m_axi_ARCACHE(m_axi_out_2_ARCACHE),
    .m_axi_ARID(m_axi_out_2_ARID),
    .m_axi_ARLEN(m_axi_out_2_ARLEN),
    .m_axi_ARLOCK(m_axi_out_2_ARLOCK),
    .m_axi_ARPROT(m_axi_out_2_ARPROT),
    .m_axi_ARQOS(m_axi_out_2_ARQOS),
    .m_axi_ARREADY(m_axi_out_2_ARREADY),
    .m_axi_ARSIZE(m_axi_out_2_ARSIZE),
    .m_axi_ARVALID(m_axi_out_2_ARVALID),
    .m_axi_AWADDR(m_axi_out_2_AWADDR),
    .m_axi_AWBURST(m_axi_out_2_AWBURST),
    .m_axi_AWCACHE(m_axi_out_2_AWCACHE),
    .m_axi_AWID(m_axi_out_2_AWID),
    .m_axi_AWLEN(m_axi_out_2_AWLEN),
    .m_axi_AWLOCK(m_axi_out_2_AWLOCK),
    .m_axi_AWPROT(m_axi_out_2_AWPROT),
    .m_axi_AWQOS(m_axi_out_2_AWQOS),
    .m_axi_AWREADY(m_axi_out_2_AWREADY),
    .m_axi_AWSIZE(m_axi_out_2_AWSIZE),
    .m_axi_AWVALID(m_axi_out_2_AWVALID),
    .m_axi_BID(m_axi_out_2_BID),
    .m_axi_BREADY(m_axi_out_2_BREADY),
    .m_axi_BRESP(m_axi_out_2_BRESP),
    .m_axi_BVALID(m_axi_out_2_BVALID),
    .m_axi_RDATA(m_axi_out_2_RDATA),
    .m_axi_RID(m_axi_out_2_RID),
    .m_axi_RLAST(m_axi_out_2_RLAST),
    .m_axi_RREADY(m_axi_out_2_RREADY),
    .m_axi_RRESP(m_axi_out_2_RRESP),
    .m_axi_RVALID(m_axi_out_2_RVALID),
    .m_axi_WDATA(m_axi_out_2_WDATA),
    .m_axi_WLAST(m_axi_out_2_WLAST),
    .m_axi_WREADY(m_axi_out_2_WREADY),
    .m_axi_WSTRB(m_axi_out_2_WSTRB),
    .m_axi_WVALID(m_axi_out_2_WVALID),
    .read_addr_din(out_2_read_addr__din),
    .read_addr_full_n(out_2_read_addr__full_n),
    .read_addr_write(out_2_read_addr__write),
    .read_data_dout(out_2_read_data__dout),
    .read_data_empty_n(out_2_read_data__empty_n),
    .read_data_read(out_2_read_data__read),
    .write_addr_din(out_2_write_addr__din),
    .write_addr_full_n(out_2_write_addr__full_n),
    .write_addr_write(out_2_write_addr__write),
    .write_data_din(out_2_write_data__din),
    .write_data_full_n(out_2_write_data__full_n),
    .write_data_write(out_2_write_data__write),
    .write_resp_dout(out_2_write_resp__dout),
    .write_resp_empty_n(out_2_write_resp__empty_n),
    .write_resp_read(out_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_3___in_3__q0),
    .m_axi_ARADDR(m_axi_in_3_ARADDR),
    .m_axi_ARBURST(m_axi_in_3_ARBURST),
    .m_axi_ARCACHE(m_axi_in_3_ARCACHE),
    .m_axi_ARID(m_axi_in_3_ARID),
    .m_axi_ARLEN(m_axi_in_3_ARLEN),
    .m_axi_ARLOCK(m_axi_in_3_ARLOCK),
    .m_axi_ARPROT(m_axi_in_3_ARPROT),
    .m_axi_ARQOS(m_axi_in_3_ARQOS),
    .m_axi_ARREADY(m_axi_in_3_ARREADY),
    .m_axi_ARSIZE(m_axi_in_3_ARSIZE),
    .m_axi_ARVALID(m_axi_in_3_ARVALID),
    .m_axi_AWADDR(m_axi_in_3_AWADDR),
    .m_axi_AWBURST(m_axi_in_3_AWBURST),
    .m_axi_AWCACHE(m_axi_in_3_AWCACHE),
    .m_axi_AWID(m_axi_in_3_AWID),
    .m_axi_AWLEN(m_axi_in_3_AWLEN),
    .m_axi_AWLOCK(m_axi_in_3_AWLOCK),
    .m_axi_AWPROT(m_axi_in_3_AWPROT),
    .m_axi_AWQOS(m_axi_in_3_AWQOS),
    .m_axi_AWREADY(m_axi_in_3_AWREADY),
    .m_axi_AWSIZE(m_axi_in_3_AWSIZE),
    .m_axi_AWVALID(m_axi_in_3_AWVALID),
    .m_axi_BID(m_axi_in_3_BID),
    .m_axi_BREADY(m_axi_in_3_BREADY),
    .m_axi_BRESP(m_axi_in_3_BRESP),
    .m_axi_BVALID(m_axi_in_3_BVALID),
    .m_axi_RDATA(m_axi_in_3_RDATA),
    .m_axi_RID(m_axi_in_3_RID),
    .m_axi_RLAST(m_axi_in_3_RLAST),
    .m_axi_RREADY(m_axi_in_3_RREADY),
    .m_axi_RRESP(m_axi_in_3_RRESP),
    .m_axi_RVALID(m_axi_in_3_RVALID),
    .m_axi_WDATA(m_axi_in_3_WDATA),
    .m_axi_WLAST(m_axi_in_3_WLAST),
    .m_axi_WREADY(m_axi_in_3_WREADY),
    .m_axi_WSTRB(m_axi_in_3_WSTRB),
    .m_axi_WVALID(m_axi_in_3_WVALID),
    .read_addr_din(in_3_read_addr__din),
    .read_addr_full_n(in_3_read_addr__full_n),
    .read_addr_write(in_3_read_addr__write),
    .read_data_dout(in_3_read_data__dout),
    .read_data_empty_n(in_3_read_data__empty_n),
    .read_data_read(in_3_read_data__read),
    .write_addr_din(in_3_write_addr__din),
    .write_addr_full_n(in_3_write_addr__full_n),
    .write_addr_write(in_3_write_addr__write),
    .write_data_din(in_3_write_data__din),
    .write_data_full_n(in_3_write_data__full_n),
    .write_data_write(in_3_write_data__write),
    .write_resp_dout(in_3_write_resp__dout),
    .write_resp_empty_n(in_3_write_resp__empty_n),
    .write_resp_read(in_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_3___out_3__q0),
    .m_axi_ARADDR(m_axi_out_3_ARADDR),
    .m_axi_ARBURST(m_axi_out_3_ARBURST),
    .m_axi_ARCACHE(m_axi_out_3_ARCACHE),
    .m_axi_ARID(m_axi_out_3_ARID),
    .m_axi_ARLEN(m_axi_out_3_ARLEN),
    .m_axi_ARLOCK(m_axi_out_3_ARLOCK),
    .m_axi_ARPROT(m_axi_out_3_ARPROT),
    .m_axi_ARQOS(m_axi_out_3_ARQOS),
    .m_axi_ARREADY(m_axi_out_3_ARREADY),
    .m_axi_ARSIZE(m_axi_out_3_ARSIZE),
    .m_axi_ARVALID(m_axi_out_3_ARVALID),
    .m_axi_AWADDR(m_axi_out_3_AWADDR),
    .m_axi_AWBURST(m_axi_out_3_AWBURST),
    .m_axi_AWCACHE(m_axi_out_3_AWCACHE),
    .m_axi_AWID(m_axi_out_3_AWID),
    .m_axi_AWLEN(m_axi_out_3_AWLEN),
    .m_axi_AWLOCK(m_axi_out_3_AWLOCK),
    .m_axi_AWPROT(m_axi_out_3_AWPROT),
    .m_axi_AWQOS(m_axi_out_3_AWQOS),
    .m_axi_AWREADY(m_axi_out_3_AWREADY),
    .m_axi_AWSIZE(m_axi_out_3_AWSIZE),
    .m_axi_AWVALID(m_axi_out_3_AWVALID),
    .m_axi_BID(m_axi_out_3_BID),
    .m_axi_BREADY(m_axi_out_3_BREADY),
    .m_axi_BRESP(m_axi_out_3_BRESP),
    .m_axi_BVALID(m_axi_out_3_BVALID),
    .m_axi_RDATA(m_axi_out_3_RDATA),
    .m_axi_RID(m_axi_out_3_RID),
    .m_axi_RLAST(m_axi_out_3_RLAST),
    .m_axi_RREADY(m_axi_out_3_RREADY),
    .m_axi_RRESP(m_axi_out_3_RRESP),
    .m_axi_RVALID(m_axi_out_3_RVALID),
    .m_axi_WDATA(m_axi_out_3_WDATA),
    .m_axi_WLAST(m_axi_out_3_WLAST),
    .m_axi_WREADY(m_axi_out_3_WREADY),
    .m_axi_WSTRB(m_axi_out_3_WSTRB),
    .m_axi_WVALID(m_axi_out_3_WVALID),
    .read_addr_din(out_3_read_addr__din),
    .read_addr_full_n(out_3_read_addr__full_n),
    .read_addr_write(out_3_read_addr__write),
    .read_data_dout(out_3_read_data__dout),
    .read_data_empty_n(out_3_read_data__empty_n),
    .read_data_read(out_3_read_data__read),
    .write_addr_din(out_3_write_addr__din),
    .write_addr_full_n(out_3_write_addr__full_n),
    .write_addr_write(out_3_write_addr__write),
    .write_data_din(out_3_write_data__din),
    .write_data_full_n(out_3_write_data__full_n),
    .write_data_write(out_3_write_data__write),
    .write_resp_dout(out_3_write_resp__dout),
    .write_resp_empty_n(out_3_write_resp__empty_n),
    .write_resp_read(out_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_4__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_4___in_4__q0),
    .m_axi_ARADDR(m_axi_in_4_ARADDR),
    .m_axi_ARBURST(m_axi_in_4_ARBURST),
    .m_axi_ARCACHE(m_axi_in_4_ARCACHE),
    .m_axi_ARID(m_axi_in_4_ARID),
    .m_axi_ARLEN(m_axi_in_4_ARLEN),
    .m_axi_ARLOCK(m_axi_in_4_ARLOCK),
    .m_axi_ARPROT(m_axi_in_4_ARPROT),
    .m_axi_ARQOS(m_axi_in_4_ARQOS),
    .m_axi_ARREADY(m_axi_in_4_ARREADY),
    .m_axi_ARSIZE(m_axi_in_4_ARSIZE),
    .m_axi_ARVALID(m_axi_in_4_ARVALID),
    .m_axi_AWADDR(m_axi_in_4_AWADDR),
    .m_axi_AWBURST(m_axi_in_4_AWBURST),
    .m_axi_AWCACHE(m_axi_in_4_AWCACHE),
    .m_axi_AWID(m_axi_in_4_AWID),
    .m_axi_AWLEN(m_axi_in_4_AWLEN),
    .m_axi_AWLOCK(m_axi_in_4_AWLOCK),
    .m_axi_AWPROT(m_axi_in_4_AWPROT),
    .m_axi_AWQOS(m_axi_in_4_AWQOS),
    .m_axi_AWREADY(m_axi_in_4_AWREADY),
    .m_axi_AWSIZE(m_axi_in_4_AWSIZE),
    .m_axi_AWVALID(m_axi_in_4_AWVALID),
    .m_axi_BID(m_axi_in_4_BID),
    .m_axi_BREADY(m_axi_in_4_BREADY),
    .m_axi_BRESP(m_axi_in_4_BRESP),
    .m_axi_BVALID(m_axi_in_4_BVALID),
    .m_axi_RDATA(m_axi_in_4_RDATA),
    .m_axi_RID(m_axi_in_4_RID),
    .m_axi_RLAST(m_axi_in_4_RLAST),
    .m_axi_RREADY(m_axi_in_4_RREADY),
    .m_axi_RRESP(m_axi_in_4_RRESP),
    .m_axi_RVALID(m_axi_in_4_RVALID),
    .m_axi_WDATA(m_axi_in_4_WDATA),
    .m_axi_WLAST(m_axi_in_4_WLAST),
    .m_axi_WREADY(m_axi_in_4_WREADY),
    .m_axi_WSTRB(m_axi_in_4_WSTRB),
    .m_axi_WVALID(m_axi_in_4_WVALID),
    .read_addr_din(in_4_read_addr__din),
    .read_addr_full_n(in_4_read_addr__full_n),
    .read_addr_write(in_4_read_addr__write),
    .read_data_dout(in_4_read_data__dout),
    .read_data_empty_n(in_4_read_data__empty_n),
    .read_data_read(in_4_read_data__read),
    .write_addr_din(in_4_write_addr__din),
    .write_addr_full_n(in_4_write_addr__full_n),
    .write_addr_write(in_4_write_addr__write),
    .write_data_din(in_4_write_data__din),
    .write_data_full_n(in_4_write_data__full_n),
    .write_data_write(in_4_write_data__write),
    .write_resp_dout(in_4_write_resp__dout),
    .write_resp_empty_n(in_4_write_resp__empty_n),
    .write_resp_read(in_4_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_4__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_4___out_4__q0),
    .m_axi_ARADDR(m_axi_out_4_ARADDR),
    .m_axi_ARBURST(m_axi_out_4_ARBURST),
    .m_axi_ARCACHE(m_axi_out_4_ARCACHE),
    .m_axi_ARID(m_axi_out_4_ARID),
    .m_axi_ARLEN(m_axi_out_4_ARLEN),
    .m_axi_ARLOCK(m_axi_out_4_ARLOCK),
    .m_axi_ARPROT(m_axi_out_4_ARPROT),
    .m_axi_ARQOS(m_axi_out_4_ARQOS),
    .m_axi_ARREADY(m_axi_out_4_ARREADY),
    .m_axi_ARSIZE(m_axi_out_4_ARSIZE),
    .m_axi_ARVALID(m_axi_out_4_ARVALID),
    .m_axi_AWADDR(m_axi_out_4_AWADDR),
    .m_axi_AWBURST(m_axi_out_4_AWBURST),
    .m_axi_AWCACHE(m_axi_out_4_AWCACHE),
    .m_axi_AWID(m_axi_out_4_AWID),
    .m_axi_AWLEN(m_axi_out_4_AWLEN),
    .m_axi_AWLOCK(m_axi_out_4_AWLOCK),
    .m_axi_AWPROT(m_axi_out_4_AWPROT),
    .m_axi_AWQOS(m_axi_out_4_AWQOS),
    .m_axi_AWREADY(m_axi_out_4_AWREADY),
    .m_axi_AWSIZE(m_axi_out_4_AWSIZE),
    .m_axi_AWVALID(m_axi_out_4_AWVALID),
    .m_axi_BID(m_axi_out_4_BID),
    .m_axi_BREADY(m_axi_out_4_BREADY),
    .m_axi_BRESP(m_axi_out_4_BRESP),
    .m_axi_BVALID(m_axi_out_4_BVALID),
    .m_axi_RDATA(m_axi_out_4_RDATA),
    .m_axi_RID(m_axi_out_4_RID),
    .m_axi_RLAST(m_axi_out_4_RLAST),
    .m_axi_RREADY(m_axi_out_4_RREADY),
    .m_axi_RRESP(m_axi_out_4_RRESP),
    .m_axi_RVALID(m_axi_out_4_RVALID),
    .m_axi_WDATA(m_axi_out_4_WDATA),
    .m_axi_WLAST(m_axi_out_4_WLAST),
    .m_axi_WREADY(m_axi_out_4_WREADY),
    .m_axi_WSTRB(m_axi_out_4_WSTRB),
    .m_axi_WVALID(m_axi_out_4_WVALID),
    .read_addr_din(out_4_read_addr__din),
    .read_addr_full_n(out_4_read_addr__full_n),
    .read_addr_write(out_4_read_addr__write),
    .read_data_dout(out_4_read_data__dout),
    .read_data_empty_n(out_4_read_data__empty_n),
    .read_data_read(out_4_read_data__read),
    .write_addr_din(out_4_write_addr__din),
    .write_addr_full_n(out_4_write_addr__full_n),
    .write_addr_write(out_4_write_addr__write),
    .write_data_din(out_4_write_data__din),
    .write_data_full_n(out_4_write_data__full_n),
    .write_data_write(out_4_write_data__write),
    .write_resp_dout(out_4_write_resp__dout),
    .write_resp_empty_n(out_4_write_resp__empty_n),
    .write_resp_read(out_4_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_5__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_5___in_5__q0),
    .m_axi_ARADDR(m_axi_in_5_ARADDR),
    .m_axi_ARBURST(m_axi_in_5_ARBURST),
    .m_axi_ARCACHE(m_axi_in_5_ARCACHE),
    .m_axi_ARID(m_axi_in_5_ARID),
    .m_axi_ARLEN(m_axi_in_5_ARLEN),
    .m_axi_ARLOCK(m_axi_in_5_ARLOCK),
    .m_axi_ARPROT(m_axi_in_5_ARPROT),
    .m_axi_ARQOS(m_axi_in_5_ARQOS),
    .m_axi_ARREADY(m_axi_in_5_ARREADY),
    .m_axi_ARSIZE(m_axi_in_5_ARSIZE),
    .m_axi_ARVALID(m_axi_in_5_ARVALID),
    .m_axi_AWADDR(m_axi_in_5_AWADDR),
    .m_axi_AWBURST(m_axi_in_5_AWBURST),
    .m_axi_AWCACHE(m_axi_in_5_AWCACHE),
    .m_axi_AWID(m_axi_in_5_AWID),
    .m_axi_AWLEN(m_axi_in_5_AWLEN),
    .m_axi_AWLOCK(m_axi_in_5_AWLOCK),
    .m_axi_AWPROT(m_axi_in_5_AWPROT),
    .m_axi_AWQOS(m_axi_in_5_AWQOS),
    .m_axi_AWREADY(m_axi_in_5_AWREADY),
    .m_axi_AWSIZE(m_axi_in_5_AWSIZE),
    .m_axi_AWVALID(m_axi_in_5_AWVALID),
    .m_axi_BID(m_axi_in_5_BID),
    .m_axi_BREADY(m_axi_in_5_BREADY),
    .m_axi_BRESP(m_axi_in_5_BRESP),
    .m_axi_BVALID(m_axi_in_5_BVALID),
    .m_axi_RDATA(m_axi_in_5_RDATA),
    .m_axi_RID(m_axi_in_5_RID),
    .m_axi_RLAST(m_axi_in_5_RLAST),
    .m_axi_RREADY(m_axi_in_5_RREADY),
    .m_axi_RRESP(m_axi_in_5_RRESP),
    .m_axi_RVALID(m_axi_in_5_RVALID),
    .m_axi_WDATA(m_axi_in_5_WDATA),
    .m_axi_WLAST(m_axi_in_5_WLAST),
    .m_axi_WREADY(m_axi_in_5_WREADY),
    .m_axi_WSTRB(m_axi_in_5_WSTRB),
    .m_axi_WVALID(m_axi_in_5_WVALID),
    .read_addr_din(in_5_read_addr__din),
    .read_addr_full_n(in_5_read_addr__full_n),
    .read_addr_write(in_5_read_addr__write),
    .read_data_dout(in_5_read_data__dout),
    .read_data_empty_n(in_5_read_data__empty_n),
    .read_data_read(in_5_read_data__read),
    .write_addr_din(in_5_write_addr__din),
    .write_addr_full_n(in_5_write_addr__full_n),
    .write_addr_write(in_5_write_addr__write),
    .write_data_din(in_5_write_data__din),
    .write_data_full_n(in_5_write_data__full_n),
    .write_data_write(in_5_write_data__write),
    .write_resp_dout(in_5_write_resp__dout),
    .write_resp_empty_n(in_5_write_resp__empty_n),
    .write_resp_read(in_5_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_5__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_5___out_5__q0),
    .m_axi_ARADDR(m_axi_out_5_ARADDR),
    .m_axi_ARBURST(m_axi_out_5_ARBURST),
    .m_axi_ARCACHE(m_axi_out_5_ARCACHE),
    .m_axi_ARID(m_axi_out_5_ARID),
    .m_axi_ARLEN(m_axi_out_5_ARLEN),
    .m_axi_ARLOCK(m_axi_out_5_ARLOCK),
    .m_axi_ARPROT(m_axi_out_5_ARPROT),
    .m_axi_ARQOS(m_axi_out_5_ARQOS),
    .m_axi_ARREADY(m_axi_out_5_ARREADY),
    .m_axi_ARSIZE(m_axi_out_5_ARSIZE),
    .m_axi_ARVALID(m_axi_out_5_ARVALID),
    .m_axi_AWADDR(m_axi_out_5_AWADDR),
    .m_axi_AWBURST(m_axi_out_5_AWBURST),
    .m_axi_AWCACHE(m_axi_out_5_AWCACHE),
    .m_axi_AWID(m_axi_out_5_AWID),
    .m_axi_AWLEN(m_axi_out_5_AWLEN),
    .m_axi_AWLOCK(m_axi_out_5_AWLOCK),
    .m_axi_AWPROT(m_axi_out_5_AWPROT),
    .m_axi_AWQOS(m_axi_out_5_AWQOS),
    .m_axi_AWREADY(m_axi_out_5_AWREADY),
    .m_axi_AWSIZE(m_axi_out_5_AWSIZE),
    .m_axi_AWVALID(m_axi_out_5_AWVALID),
    .m_axi_BID(m_axi_out_5_BID),
    .m_axi_BREADY(m_axi_out_5_BREADY),
    .m_axi_BRESP(m_axi_out_5_BRESP),
    .m_axi_BVALID(m_axi_out_5_BVALID),
    .m_axi_RDATA(m_axi_out_5_RDATA),
    .m_axi_RID(m_axi_out_5_RID),
    .m_axi_RLAST(m_axi_out_5_RLAST),
    .m_axi_RREADY(m_axi_out_5_RREADY),
    .m_axi_RRESP(m_axi_out_5_RRESP),
    .m_axi_RVALID(m_axi_out_5_RVALID),
    .m_axi_WDATA(m_axi_out_5_WDATA),
    .m_axi_WLAST(m_axi_out_5_WLAST),
    .m_axi_WREADY(m_axi_out_5_WREADY),
    .m_axi_WSTRB(m_axi_out_5_WSTRB),
    .m_axi_WVALID(m_axi_out_5_WVALID),
    .read_addr_din(out_5_read_addr__din),
    .read_addr_full_n(out_5_read_addr__full_n),
    .read_addr_write(out_5_read_addr__write),
    .read_data_dout(out_5_read_data__dout),
    .read_data_empty_n(out_5_read_data__empty_n),
    .read_data_read(out_5_read_data__read),
    .write_addr_din(out_5_write_addr__din),
    .write_addr_full_n(out_5_write_addr__full_n),
    .write_addr_write(out_5_write_addr__write),
    .write_data_din(out_5_write_data__din),
    .write_data_full_n(out_5_write_data__full_n),
    .write_data_write(out_5_write_data__write),
    .write_resp_dout(out_5_write_resp__dout),
    .write_resp_empty_n(out_5_write_resp__empty_n),
    .write_resp_read(out_5_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_6__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_6___in_6__q0),
    .m_axi_ARADDR(m_axi_in_6_ARADDR),
    .m_axi_ARBURST(m_axi_in_6_ARBURST),
    .m_axi_ARCACHE(m_axi_in_6_ARCACHE),
    .m_axi_ARID(m_axi_in_6_ARID),
    .m_axi_ARLEN(m_axi_in_6_ARLEN),
    .m_axi_ARLOCK(m_axi_in_6_ARLOCK),
    .m_axi_ARPROT(m_axi_in_6_ARPROT),
    .m_axi_ARQOS(m_axi_in_6_ARQOS),
    .m_axi_ARREADY(m_axi_in_6_ARREADY),
    .m_axi_ARSIZE(m_axi_in_6_ARSIZE),
    .m_axi_ARVALID(m_axi_in_6_ARVALID),
    .m_axi_AWADDR(m_axi_in_6_AWADDR),
    .m_axi_AWBURST(m_axi_in_6_AWBURST),
    .m_axi_AWCACHE(m_axi_in_6_AWCACHE),
    .m_axi_AWID(m_axi_in_6_AWID),
    .m_axi_AWLEN(m_axi_in_6_AWLEN),
    .m_axi_AWLOCK(m_axi_in_6_AWLOCK),
    .m_axi_AWPROT(m_axi_in_6_AWPROT),
    .m_axi_AWQOS(m_axi_in_6_AWQOS),
    .m_axi_AWREADY(m_axi_in_6_AWREADY),
    .m_axi_AWSIZE(m_axi_in_6_AWSIZE),
    .m_axi_AWVALID(m_axi_in_6_AWVALID),
    .m_axi_BID(m_axi_in_6_BID),
    .m_axi_BREADY(m_axi_in_6_BREADY),
    .m_axi_BRESP(m_axi_in_6_BRESP),
    .m_axi_BVALID(m_axi_in_6_BVALID),
    .m_axi_RDATA(m_axi_in_6_RDATA),
    .m_axi_RID(m_axi_in_6_RID),
    .m_axi_RLAST(m_axi_in_6_RLAST),
    .m_axi_RREADY(m_axi_in_6_RREADY),
    .m_axi_RRESP(m_axi_in_6_RRESP),
    .m_axi_RVALID(m_axi_in_6_RVALID),
    .m_axi_WDATA(m_axi_in_6_WDATA),
    .m_axi_WLAST(m_axi_in_6_WLAST),
    .m_axi_WREADY(m_axi_in_6_WREADY),
    .m_axi_WSTRB(m_axi_in_6_WSTRB),
    .m_axi_WVALID(m_axi_in_6_WVALID),
    .read_addr_din(in_6_read_addr__din),
    .read_addr_full_n(in_6_read_addr__full_n),
    .read_addr_write(in_6_read_addr__write),
    .read_data_dout(in_6_read_data__dout),
    .read_data_empty_n(in_6_read_data__empty_n),
    .read_data_read(in_6_read_data__read),
    .write_addr_din(in_6_write_addr__din),
    .write_addr_full_n(in_6_write_addr__full_n),
    .write_addr_write(in_6_write_addr__write),
    .write_data_din(in_6_write_data__din),
    .write_data_full_n(in_6_write_data__full_n),
    .write_data_write(in_6_write_data__write),
    .write_resp_dout(in_6_write_resp__dout),
    .write_resp_empty_n(in_6_write_resp__empty_n),
    .write_resp_read(in_6_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_6__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_6___out_6__q0),
    .m_axi_ARADDR(m_axi_out_6_ARADDR),
    .m_axi_ARBURST(m_axi_out_6_ARBURST),
    .m_axi_ARCACHE(m_axi_out_6_ARCACHE),
    .m_axi_ARID(m_axi_out_6_ARID),
    .m_axi_ARLEN(m_axi_out_6_ARLEN),
    .m_axi_ARLOCK(m_axi_out_6_ARLOCK),
    .m_axi_ARPROT(m_axi_out_6_ARPROT),
    .m_axi_ARQOS(m_axi_out_6_ARQOS),
    .m_axi_ARREADY(m_axi_out_6_ARREADY),
    .m_axi_ARSIZE(m_axi_out_6_ARSIZE),
    .m_axi_ARVALID(m_axi_out_6_ARVALID),
    .m_axi_AWADDR(m_axi_out_6_AWADDR),
    .m_axi_AWBURST(m_axi_out_6_AWBURST),
    .m_axi_AWCACHE(m_axi_out_6_AWCACHE),
    .m_axi_AWID(m_axi_out_6_AWID),
    .m_axi_AWLEN(m_axi_out_6_AWLEN),
    .m_axi_AWLOCK(m_axi_out_6_AWLOCK),
    .m_axi_AWPROT(m_axi_out_6_AWPROT),
    .m_axi_AWQOS(m_axi_out_6_AWQOS),
    .m_axi_AWREADY(m_axi_out_6_AWREADY),
    .m_axi_AWSIZE(m_axi_out_6_AWSIZE),
    .m_axi_AWVALID(m_axi_out_6_AWVALID),
    .m_axi_BID(m_axi_out_6_BID),
    .m_axi_BREADY(m_axi_out_6_BREADY),
    .m_axi_BRESP(m_axi_out_6_BRESP),
    .m_axi_BVALID(m_axi_out_6_BVALID),
    .m_axi_RDATA(m_axi_out_6_RDATA),
    .m_axi_RID(m_axi_out_6_RID),
    .m_axi_RLAST(m_axi_out_6_RLAST),
    .m_axi_RREADY(m_axi_out_6_RREADY),
    .m_axi_RRESP(m_axi_out_6_RRESP),
    .m_axi_RVALID(m_axi_out_6_RVALID),
    .m_axi_WDATA(m_axi_out_6_WDATA),
    .m_axi_WLAST(m_axi_out_6_WLAST),
    .m_axi_WREADY(m_axi_out_6_WREADY),
    .m_axi_WSTRB(m_axi_out_6_WSTRB),
    .m_axi_WVALID(m_axi_out_6_WVALID),
    .read_addr_din(out_6_read_addr__din),
    .read_addr_full_n(out_6_read_addr__full_n),
    .read_addr_write(out_6_read_addr__write),
    .read_data_dout(out_6_read_data__dout),
    .read_data_empty_n(out_6_read_data__empty_n),
    .read_data_read(out_6_read_data__read),
    .write_addr_din(out_6_write_addr__din),
    .write_addr_full_n(out_6_write_addr__full_n),
    .write_addr_write(out_6_write_addr__write),
    .write_data_din(out_6_write_data__din),
    .write_data_full_n(out_6_write_data__full_n),
    .write_data_write(out_6_write_data__write),
    .write_resp_dout(out_6_write_resp__dout),
    .write_resp_empty_n(out_6_write_resp__empty_n),
    .write_resp_read(out_6_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_7__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_7___in_7__q0),
    .m_axi_ARADDR(m_axi_in_7_ARADDR),
    .m_axi_ARBURST(m_axi_in_7_ARBURST),
    .m_axi_ARCACHE(m_axi_in_7_ARCACHE),
    .m_axi_ARID(m_axi_in_7_ARID),
    .m_axi_ARLEN(m_axi_in_7_ARLEN),
    .m_axi_ARLOCK(m_axi_in_7_ARLOCK),
    .m_axi_ARPROT(m_axi_in_7_ARPROT),
    .m_axi_ARQOS(m_axi_in_7_ARQOS),
    .m_axi_ARREADY(m_axi_in_7_ARREADY),
    .m_axi_ARSIZE(m_axi_in_7_ARSIZE),
    .m_axi_ARVALID(m_axi_in_7_ARVALID),
    .m_axi_AWADDR(m_axi_in_7_AWADDR),
    .m_axi_AWBURST(m_axi_in_7_AWBURST),
    .m_axi_AWCACHE(m_axi_in_7_AWCACHE),
    .m_axi_AWID(m_axi_in_7_AWID),
    .m_axi_AWLEN(m_axi_in_7_AWLEN),
    .m_axi_AWLOCK(m_axi_in_7_AWLOCK),
    .m_axi_AWPROT(m_axi_in_7_AWPROT),
    .m_axi_AWQOS(m_axi_in_7_AWQOS),
    .m_axi_AWREADY(m_axi_in_7_AWREADY),
    .m_axi_AWSIZE(m_axi_in_7_AWSIZE),
    .m_axi_AWVALID(m_axi_in_7_AWVALID),
    .m_axi_BID(m_axi_in_7_BID),
    .m_axi_BREADY(m_axi_in_7_BREADY),
    .m_axi_BRESP(m_axi_in_7_BRESP),
    .m_axi_BVALID(m_axi_in_7_BVALID),
    .m_axi_RDATA(m_axi_in_7_RDATA),
    .m_axi_RID(m_axi_in_7_RID),
    .m_axi_RLAST(m_axi_in_7_RLAST),
    .m_axi_RREADY(m_axi_in_7_RREADY),
    .m_axi_RRESP(m_axi_in_7_RRESP),
    .m_axi_RVALID(m_axi_in_7_RVALID),
    .m_axi_WDATA(m_axi_in_7_WDATA),
    .m_axi_WLAST(m_axi_in_7_WLAST),
    .m_axi_WREADY(m_axi_in_7_WREADY),
    .m_axi_WSTRB(m_axi_in_7_WSTRB),
    .m_axi_WVALID(m_axi_in_7_WVALID),
    .read_addr_din(in_7_read_addr__din),
    .read_addr_full_n(in_7_read_addr__full_n),
    .read_addr_write(in_7_read_addr__write),
    .read_data_dout(in_7_read_data__dout),
    .read_data_empty_n(in_7_read_data__empty_n),
    .read_data_read(in_7_read_data__read),
    .write_addr_din(in_7_write_addr__din),
    .write_addr_full_n(in_7_write_addr__full_n),
    .write_addr_write(in_7_write_addr__write),
    .write_data_din(in_7_write_data__din),
    .write_data_full_n(in_7_write_data__full_n),
    .write_data_write(in_7_write_data__write),
    .write_resp_dout(in_7_write_resp__dout),
    .write_resp_empty_n(in_7_write_resp__empty_n),
    .write_resp_read(in_7_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_7__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_7___out_7__q0),
    .m_axi_ARADDR(m_axi_out_7_ARADDR),
    .m_axi_ARBURST(m_axi_out_7_ARBURST),
    .m_axi_ARCACHE(m_axi_out_7_ARCACHE),
    .m_axi_ARID(m_axi_out_7_ARID),
    .m_axi_ARLEN(m_axi_out_7_ARLEN),
    .m_axi_ARLOCK(m_axi_out_7_ARLOCK),
    .m_axi_ARPROT(m_axi_out_7_ARPROT),
    .m_axi_ARQOS(m_axi_out_7_ARQOS),
    .m_axi_ARREADY(m_axi_out_7_ARREADY),
    .m_axi_ARSIZE(m_axi_out_7_ARSIZE),
    .m_axi_ARVALID(m_axi_out_7_ARVALID),
    .m_axi_AWADDR(m_axi_out_7_AWADDR),
    .m_axi_AWBURST(m_axi_out_7_AWBURST),
    .m_axi_AWCACHE(m_axi_out_7_AWCACHE),
    .m_axi_AWID(m_axi_out_7_AWID),
    .m_axi_AWLEN(m_axi_out_7_AWLEN),
    .m_axi_AWLOCK(m_axi_out_7_AWLOCK),
    .m_axi_AWPROT(m_axi_out_7_AWPROT),
    .m_axi_AWQOS(m_axi_out_7_AWQOS),
    .m_axi_AWREADY(m_axi_out_7_AWREADY),
    .m_axi_AWSIZE(m_axi_out_7_AWSIZE),
    .m_axi_AWVALID(m_axi_out_7_AWVALID),
    .m_axi_BID(m_axi_out_7_BID),
    .m_axi_BREADY(m_axi_out_7_BREADY),
    .m_axi_BRESP(m_axi_out_7_BRESP),
    .m_axi_BVALID(m_axi_out_7_BVALID),
    .m_axi_RDATA(m_axi_out_7_RDATA),
    .m_axi_RID(m_axi_out_7_RID),
    .m_axi_RLAST(m_axi_out_7_RLAST),
    .m_axi_RREADY(m_axi_out_7_RREADY),
    .m_axi_RRESP(m_axi_out_7_RRESP),
    .m_axi_RVALID(m_axi_out_7_RVALID),
    .m_axi_WDATA(m_axi_out_7_WDATA),
    .m_axi_WLAST(m_axi_out_7_WLAST),
    .m_axi_WREADY(m_axi_out_7_WREADY),
    .m_axi_WSTRB(m_axi_out_7_WSTRB),
    .m_axi_WVALID(m_axi_out_7_WVALID),
    .read_addr_din(out_7_read_addr__din),
    .read_addr_full_n(out_7_read_addr__full_n),
    .read_addr_write(out_7_read_addr__write),
    .read_data_dout(out_7_read_data__dout),
    .read_data_empty_n(out_7_read_data__empty_n),
    .read_data_read(out_7_read_data__read),
    .write_addr_din(out_7_write_addr__din),
    .write_addr_full_n(out_7_write_addr__full_n),
    .write_addr_write(out_7_write_addr__write),
    .write_data_din(out_7_write_data__din),
    .write_data_full_n(out_7_write_data__full_n),
    .write_data_write(out_7_write_data__write),
    .write_resp_dout(out_7_write_resp__dout),
    .write_resp_empty_n(out_7_write_resp__empty_n),
    .write_resp_read(out_7_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_8__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_8___in_8__q0),
    .m_axi_ARADDR(m_axi_in_8_ARADDR),
    .m_axi_ARBURST(m_axi_in_8_ARBURST),
    .m_axi_ARCACHE(m_axi_in_8_ARCACHE),
    .m_axi_ARID(m_axi_in_8_ARID),
    .m_axi_ARLEN(m_axi_in_8_ARLEN),
    .m_axi_ARLOCK(m_axi_in_8_ARLOCK),
    .m_axi_ARPROT(m_axi_in_8_ARPROT),
    .m_axi_ARQOS(m_axi_in_8_ARQOS),
    .m_axi_ARREADY(m_axi_in_8_ARREADY),
    .m_axi_ARSIZE(m_axi_in_8_ARSIZE),
    .m_axi_ARVALID(m_axi_in_8_ARVALID),
    .m_axi_AWADDR(m_axi_in_8_AWADDR),
    .m_axi_AWBURST(m_axi_in_8_AWBURST),
    .m_axi_AWCACHE(m_axi_in_8_AWCACHE),
    .m_axi_AWID(m_axi_in_8_AWID),
    .m_axi_AWLEN(m_axi_in_8_AWLEN),
    .m_axi_AWLOCK(m_axi_in_8_AWLOCK),
    .m_axi_AWPROT(m_axi_in_8_AWPROT),
    .m_axi_AWQOS(m_axi_in_8_AWQOS),
    .m_axi_AWREADY(m_axi_in_8_AWREADY),
    .m_axi_AWSIZE(m_axi_in_8_AWSIZE),
    .m_axi_AWVALID(m_axi_in_8_AWVALID),
    .m_axi_BID(m_axi_in_8_BID),
    .m_axi_BREADY(m_axi_in_8_BREADY),
    .m_axi_BRESP(m_axi_in_8_BRESP),
    .m_axi_BVALID(m_axi_in_8_BVALID),
    .m_axi_RDATA(m_axi_in_8_RDATA),
    .m_axi_RID(m_axi_in_8_RID),
    .m_axi_RLAST(m_axi_in_8_RLAST),
    .m_axi_RREADY(m_axi_in_8_RREADY),
    .m_axi_RRESP(m_axi_in_8_RRESP),
    .m_axi_RVALID(m_axi_in_8_RVALID),
    .m_axi_WDATA(m_axi_in_8_WDATA),
    .m_axi_WLAST(m_axi_in_8_WLAST),
    .m_axi_WREADY(m_axi_in_8_WREADY),
    .m_axi_WSTRB(m_axi_in_8_WSTRB),
    .m_axi_WVALID(m_axi_in_8_WVALID),
    .read_addr_din(in_8_read_addr__din),
    .read_addr_full_n(in_8_read_addr__full_n),
    .read_addr_write(in_8_read_addr__write),
    .read_data_dout(in_8_read_data__dout),
    .read_data_empty_n(in_8_read_data__empty_n),
    .read_data_read(in_8_read_data__read),
    .write_addr_din(in_8_write_addr__din),
    .write_addr_full_n(in_8_write_addr__full_n),
    .write_addr_write(in_8_write_addr__write),
    .write_data_din(in_8_write_data__din),
    .write_data_full_n(in_8_write_data__full_n),
    .write_data_write(in_8_write_data__write),
    .write_resp_dout(in_8_write_resp__dout),
    .write_resp_empty_n(in_8_write_resp__empty_n),
    .write_resp_read(in_8_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_8__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_8___out_8__q0),
    .m_axi_ARADDR(m_axi_out_8_ARADDR),
    .m_axi_ARBURST(m_axi_out_8_ARBURST),
    .m_axi_ARCACHE(m_axi_out_8_ARCACHE),
    .m_axi_ARID(m_axi_out_8_ARID),
    .m_axi_ARLEN(m_axi_out_8_ARLEN),
    .m_axi_ARLOCK(m_axi_out_8_ARLOCK),
    .m_axi_ARPROT(m_axi_out_8_ARPROT),
    .m_axi_ARQOS(m_axi_out_8_ARQOS),
    .m_axi_ARREADY(m_axi_out_8_ARREADY),
    .m_axi_ARSIZE(m_axi_out_8_ARSIZE),
    .m_axi_ARVALID(m_axi_out_8_ARVALID),
    .m_axi_AWADDR(m_axi_out_8_AWADDR),
    .m_axi_AWBURST(m_axi_out_8_AWBURST),
    .m_axi_AWCACHE(m_axi_out_8_AWCACHE),
    .m_axi_AWID(m_axi_out_8_AWID),
    .m_axi_AWLEN(m_axi_out_8_AWLEN),
    .m_axi_AWLOCK(m_axi_out_8_AWLOCK),
    .m_axi_AWPROT(m_axi_out_8_AWPROT),
    .m_axi_AWQOS(m_axi_out_8_AWQOS),
    .m_axi_AWREADY(m_axi_out_8_AWREADY),
    .m_axi_AWSIZE(m_axi_out_8_AWSIZE),
    .m_axi_AWVALID(m_axi_out_8_AWVALID),
    .m_axi_BID(m_axi_out_8_BID),
    .m_axi_BREADY(m_axi_out_8_BREADY),
    .m_axi_BRESP(m_axi_out_8_BRESP),
    .m_axi_BVALID(m_axi_out_8_BVALID),
    .m_axi_RDATA(m_axi_out_8_RDATA),
    .m_axi_RID(m_axi_out_8_RID),
    .m_axi_RLAST(m_axi_out_8_RLAST),
    .m_axi_RREADY(m_axi_out_8_RREADY),
    .m_axi_RRESP(m_axi_out_8_RRESP),
    .m_axi_RVALID(m_axi_out_8_RVALID),
    .m_axi_WDATA(m_axi_out_8_WDATA),
    .m_axi_WLAST(m_axi_out_8_WLAST),
    .m_axi_WREADY(m_axi_out_8_WREADY),
    .m_axi_WSTRB(m_axi_out_8_WSTRB),
    .m_axi_WVALID(m_axi_out_8_WVALID),
    .read_addr_din(out_8_read_addr__din),
    .read_addr_full_n(out_8_read_addr__full_n),
    .read_addr_write(out_8_read_addr__write),
    .read_data_dout(out_8_read_data__dout),
    .read_data_empty_n(out_8_read_data__empty_n),
    .read_data_read(out_8_read_data__read),
    .write_addr_din(out_8_write_addr__din),
    .write_addr_full_n(out_8_write_addr__full_n),
    .write_addr_write(out_8_write_addr__write),
    .write_data_din(out_8_write_data__din),
    .write_data_full_n(out_8_write_data__full_n),
    .write_data_write(out_8_write_data__write),
    .write_resp_dout(out_8_write_resp__dout),
    .write_resp_empty_n(out_8_write_resp__empty_n),
    .write_resp_read(out_8_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_9__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_9___in_9__q0),
    .m_axi_ARADDR(m_axi_in_9_ARADDR),
    .m_axi_ARBURST(m_axi_in_9_ARBURST),
    .m_axi_ARCACHE(m_axi_in_9_ARCACHE),
    .m_axi_ARID(m_axi_in_9_ARID),
    .m_axi_ARLEN(m_axi_in_9_ARLEN),
    .m_axi_ARLOCK(m_axi_in_9_ARLOCK),
    .m_axi_ARPROT(m_axi_in_9_ARPROT),
    .m_axi_ARQOS(m_axi_in_9_ARQOS),
    .m_axi_ARREADY(m_axi_in_9_ARREADY),
    .m_axi_ARSIZE(m_axi_in_9_ARSIZE),
    .m_axi_ARVALID(m_axi_in_9_ARVALID),
    .m_axi_AWADDR(m_axi_in_9_AWADDR),
    .m_axi_AWBURST(m_axi_in_9_AWBURST),
    .m_axi_AWCACHE(m_axi_in_9_AWCACHE),
    .m_axi_AWID(m_axi_in_9_AWID),
    .m_axi_AWLEN(m_axi_in_9_AWLEN),
    .m_axi_AWLOCK(m_axi_in_9_AWLOCK),
    .m_axi_AWPROT(m_axi_in_9_AWPROT),
    .m_axi_AWQOS(m_axi_in_9_AWQOS),
    .m_axi_AWREADY(m_axi_in_9_AWREADY),
    .m_axi_AWSIZE(m_axi_in_9_AWSIZE),
    .m_axi_AWVALID(m_axi_in_9_AWVALID),
    .m_axi_BID(m_axi_in_9_BID),
    .m_axi_BREADY(m_axi_in_9_BREADY),
    .m_axi_BRESP(m_axi_in_9_BRESP),
    .m_axi_BVALID(m_axi_in_9_BVALID),
    .m_axi_RDATA(m_axi_in_9_RDATA),
    .m_axi_RID(m_axi_in_9_RID),
    .m_axi_RLAST(m_axi_in_9_RLAST),
    .m_axi_RREADY(m_axi_in_9_RREADY),
    .m_axi_RRESP(m_axi_in_9_RRESP),
    .m_axi_RVALID(m_axi_in_9_RVALID),
    .m_axi_WDATA(m_axi_in_9_WDATA),
    .m_axi_WLAST(m_axi_in_9_WLAST),
    .m_axi_WREADY(m_axi_in_9_WREADY),
    .m_axi_WSTRB(m_axi_in_9_WSTRB),
    .m_axi_WVALID(m_axi_in_9_WVALID),
    .read_addr_din(in_9_read_addr__din),
    .read_addr_full_n(in_9_read_addr__full_n),
    .read_addr_write(in_9_read_addr__write),
    .read_data_dout(in_9_read_data__dout),
    .read_data_empty_n(in_9_read_data__empty_n),
    .read_data_read(in_9_read_data__read),
    .write_addr_din(in_9_write_addr__din),
    .write_addr_full_n(in_9_write_addr__full_n),
    .write_addr_write(in_9_write_addr__write),
    .write_data_din(in_9_write_data__din),
    .write_data_full_n(in_9_write_data__full_n),
    .write_data_write(in_9_write_data__write),
    .write_resp_dout(in_9_write_resp__dout),
    .write_resp_empty_n(in_9_write_resp__empty_n),
    .write_resp_read(in_9_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_9__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_9___out_9__q0),
    .m_axi_ARADDR(m_axi_out_9_ARADDR),
    .m_axi_ARBURST(m_axi_out_9_ARBURST),
    .m_axi_ARCACHE(m_axi_out_9_ARCACHE),
    .m_axi_ARID(m_axi_out_9_ARID),
    .m_axi_ARLEN(m_axi_out_9_ARLEN),
    .m_axi_ARLOCK(m_axi_out_9_ARLOCK),
    .m_axi_ARPROT(m_axi_out_9_ARPROT),
    .m_axi_ARQOS(m_axi_out_9_ARQOS),
    .m_axi_ARREADY(m_axi_out_9_ARREADY),
    .m_axi_ARSIZE(m_axi_out_9_ARSIZE),
    .m_axi_ARVALID(m_axi_out_9_ARVALID),
    .m_axi_AWADDR(m_axi_out_9_AWADDR),
    .m_axi_AWBURST(m_axi_out_9_AWBURST),
    .m_axi_AWCACHE(m_axi_out_9_AWCACHE),
    .m_axi_AWID(m_axi_out_9_AWID),
    .m_axi_AWLEN(m_axi_out_9_AWLEN),
    .m_axi_AWLOCK(m_axi_out_9_AWLOCK),
    .m_axi_AWPROT(m_axi_out_9_AWPROT),
    .m_axi_AWQOS(m_axi_out_9_AWQOS),
    .m_axi_AWREADY(m_axi_out_9_AWREADY),
    .m_axi_AWSIZE(m_axi_out_9_AWSIZE),
    .m_axi_AWVALID(m_axi_out_9_AWVALID),
    .m_axi_BID(m_axi_out_9_BID),
    .m_axi_BREADY(m_axi_out_9_BREADY),
    .m_axi_BRESP(m_axi_out_9_BRESP),
    .m_axi_BVALID(m_axi_out_9_BVALID),
    .m_axi_RDATA(m_axi_out_9_RDATA),
    .m_axi_RID(m_axi_out_9_RID),
    .m_axi_RLAST(m_axi_out_9_RLAST),
    .m_axi_RREADY(m_axi_out_9_RREADY),
    .m_axi_RRESP(m_axi_out_9_RRESP),
    .m_axi_RVALID(m_axi_out_9_RVALID),
    .m_axi_WDATA(m_axi_out_9_WDATA),
    .m_axi_WLAST(m_axi_out_9_WLAST),
    .m_axi_WREADY(m_axi_out_9_WREADY),
    .m_axi_WSTRB(m_axi_out_9_WSTRB),
    .m_axi_WVALID(m_axi_out_9_WVALID),
    .read_addr_din(out_9_read_addr__din),
    .read_addr_full_n(out_9_read_addr__full_n),
    .read_addr_write(out_9_read_addr__write),
    .read_data_dout(out_9_read_data__dout),
    .read_data_empty_n(out_9_read_data__empty_n),
    .read_data_read(out_9_read_data__read),
    .write_addr_din(out_9_write_addr__din),
    .write_addr_full_n(out_9_write_addr__full_n),
    .write_addr_write(out_9_write_addr__write),
    .write_data_din(out_9_write_data__din),
    .write_data_full_n(out_9_write_data__full_n),
    .write_data_write(out_9_write_data__write),
    .write_resp_dout(out_9_write_resp__dout),
    .write_resp_empty_n(out_9_write_resp__empty_n),
    .write_resp_read(out_9_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_10__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_10___in_10__q0),
    .m_axi_ARADDR(m_axi_in_10_ARADDR),
    .m_axi_ARBURST(m_axi_in_10_ARBURST),
    .m_axi_ARCACHE(m_axi_in_10_ARCACHE),
    .m_axi_ARID(m_axi_in_10_ARID),
    .m_axi_ARLEN(m_axi_in_10_ARLEN),
    .m_axi_ARLOCK(m_axi_in_10_ARLOCK),
    .m_axi_ARPROT(m_axi_in_10_ARPROT),
    .m_axi_ARQOS(m_axi_in_10_ARQOS),
    .m_axi_ARREADY(m_axi_in_10_ARREADY),
    .m_axi_ARSIZE(m_axi_in_10_ARSIZE),
    .m_axi_ARVALID(m_axi_in_10_ARVALID),
    .m_axi_AWADDR(m_axi_in_10_AWADDR),
    .m_axi_AWBURST(m_axi_in_10_AWBURST),
    .m_axi_AWCACHE(m_axi_in_10_AWCACHE),
    .m_axi_AWID(m_axi_in_10_AWID),
    .m_axi_AWLEN(m_axi_in_10_AWLEN),
    .m_axi_AWLOCK(m_axi_in_10_AWLOCK),
    .m_axi_AWPROT(m_axi_in_10_AWPROT),
    .m_axi_AWQOS(m_axi_in_10_AWQOS),
    .m_axi_AWREADY(m_axi_in_10_AWREADY),
    .m_axi_AWSIZE(m_axi_in_10_AWSIZE),
    .m_axi_AWVALID(m_axi_in_10_AWVALID),
    .m_axi_BID(m_axi_in_10_BID),
    .m_axi_BREADY(m_axi_in_10_BREADY),
    .m_axi_BRESP(m_axi_in_10_BRESP),
    .m_axi_BVALID(m_axi_in_10_BVALID),
    .m_axi_RDATA(m_axi_in_10_RDATA),
    .m_axi_RID(m_axi_in_10_RID),
    .m_axi_RLAST(m_axi_in_10_RLAST),
    .m_axi_RREADY(m_axi_in_10_RREADY),
    .m_axi_RRESP(m_axi_in_10_RRESP),
    .m_axi_RVALID(m_axi_in_10_RVALID),
    .m_axi_WDATA(m_axi_in_10_WDATA),
    .m_axi_WLAST(m_axi_in_10_WLAST),
    .m_axi_WREADY(m_axi_in_10_WREADY),
    .m_axi_WSTRB(m_axi_in_10_WSTRB),
    .m_axi_WVALID(m_axi_in_10_WVALID),
    .read_addr_din(in_10_read_addr__din),
    .read_addr_full_n(in_10_read_addr__full_n),
    .read_addr_write(in_10_read_addr__write),
    .read_data_dout(in_10_read_data__dout),
    .read_data_empty_n(in_10_read_data__empty_n),
    .read_data_read(in_10_read_data__read),
    .write_addr_din(in_10_write_addr__din),
    .write_addr_full_n(in_10_write_addr__full_n),
    .write_addr_write(in_10_write_addr__write),
    .write_data_din(in_10_write_data__din),
    .write_data_full_n(in_10_write_data__full_n),
    .write_data_write(in_10_write_data__write),
    .write_resp_dout(in_10_write_resp__dout),
    .write_resp_empty_n(in_10_write_resp__empty_n),
    .write_resp_read(in_10_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_10__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_10___out_10__q0),
    .m_axi_ARADDR(m_axi_out_10_ARADDR),
    .m_axi_ARBURST(m_axi_out_10_ARBURST),
    .m_axi_ARCACHE(m_axi_out_10_ARCACHE),
    .m_axi_ARID(m_axi_out_10_ARID),
    .m_axi_ARLEN(m_axi_out_10_ARLEN),
    .m_axi_ARLOCK(m_axi_out_10_ARLOCK),
    .m_axi_ARPROT(m_axi_out_10_ARPROT),
    .m_axi_ARQOS(m_axi_out_10_ARQOS),
    .m_axi_ARREADY(m_axi_out_10_ARREADY),
    .m_axi_ARSIZE(m_axi_out_10_ARSIZE),
    .m_axi_ARVALID(m_axi_out_10_ARVALID),
    .m_axi_AWADDR(m_axi_out_10_AWADDR),
    .m_axi_AWBURST(m_axi_out_10_AWBURST),
    .m_axi_AWCACHE(m_axi_out_10_AWCACHE),
    .m_axi_AWID(m_axi_out_10_AWID),
    .m_axi_AWLEN(m_axi_out_10_AWLEN),
    .m_axi_AWLOCK(m_axi_out_10_AWLOCK),
    .m_axi_AWPROT(m_axi_out_10_AWPROT),
    .m_axi_AWQOS(m_axi_out_10_AWQOS),
    .m_axi_AWREADY(m_axi_out_10_AWREADY),
    .m_axi_AWSIZE(m_axi_out_10_AWSIZE),
    .m_axi_AWVALID(m_axi_out_10_AWVALID),
    .m_axi_BID(m_axi_out_10_BID),
    .m_axi_BREADY(m_axi_out_10_BREADY),
    .m_axi_BRESP(m_axi_out_10_BRESP),
    .m_axi_BVALID(m_axi_out_10_BVALID),
    .m_axi_RDATA(m_axi_out_10_RDATA),
    .m_axi_RID(m_axi_out_10_RID),
    .m_axi_RLAST(m_axi_out_10_RLAST),
    .m_axi_RREADY(m_axi_out_10_RREADY),
    .m_axi_RRESP(m_axi_out_10_RRESP),
    .m_axi_RVALID(m_axi_out_10_RVALID),
    .m_axi_WDATA(m_axi_out_10_WDATA),
    .m_axi_WLAST(m_axi_out_10_WLAST),
    .m_axi_WREADY(m_axi_out_10_WREADY),
    .m_axi_WSTRB(m_axi_out_10_WSTRB),
    .m_axi_WVALID(m_axi_out_10_WVALID),
    .read_addr_din(out_10_read_addr__din),
    .read_addr_full_n(out_10_read_addr__full_n),
    .read_addr_write(out_10_read_addr__write),
    .read_data_dout(out_10_read_data__dout),
    .read_data_empty_n(out_10_read_data__empty_n),
    .read_data_read(out_10_read_data__read),
    .write_addr_din(out_10_write_addr__din),
    .write_addr_full_n(out_10_write_addr__full_n),
    .write_addr_write(out_10_write_addr__write),
    .write_data_din(out_10_write_data__din),
    .write_data_full_n(out_10_write_data__full_n),
    .write_data_write(out_10_write_data__write),
    .write_resp_dout(out_10_write_resp__dout),
    .write_resp_empty_n(out_10_write_resp__empty_n),
    .write_resp_read(out_10_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_11__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_11___in_11__q0),
    .m_axi_ARADDR(m_axi_in_11_ARADDR),
    .m_axi_ARBURST(m_axi_in_11_ARBURST),
    .m_axi_ARCACHE(m_axi_in_11_ARCACHE),
    .m_axi_ARID(m_axi_in_11_ARID),
    .m_axi_ARLEN(m_axi_in_11_ARLEN),
    .m_axi_ARLOCK(m_axi_in_11_ARLOCK),
    .m_axi_ARPROT(m_axi_in_11_ARPROT),
    .m_axi_ARQOS(m_axi_in_11_ARQOS),
    .m_axi_ARREADY(m_axi_in_11_ARREADY),
    .m_axi_ARSIZE(m_axi_in_11_ARSIZE),
    .m_axi_ARVALID(m_axi_in_11_ARVALID),
    .m_axi_AWADDR(m_axi_in_11_AWADDR),
    .m_axi_AWBURST(m_axi_in_11_AWBURST),
    .m_axi_AWCACHE(m_axi_in_11_AWCACHE),
    .m_axi_AWID(m_axi_in_11_AWID),
    .m_axi_AWLEN(m_axi_in_11_AWLEN),
    .m_axi_AWLOCK(m_axi_in_11_AWLOCK),
    .m_axi_AWPROT(m_axi_in_11_AWPROT),
    .m_axi_AWQOS(m_axi_in_11_AWQOS),
    .m_axi_AWREADY(m_axi_in_11_AWREADY),
    .m_axi_AWSIZE(m_axi_in_11_AWSIZE),
    .m_axi_AWVALID(m_axi_in_11_AWVALID),
    .m_axi_BID(m_axi_in_11_BID),
    .m_axi_BREADY(m_axi_in_11_BREADY),
    .m_axi_BRESP(m_axi_in_11_BRESP),
    .m_axi_BVALID(m_axi_in_11_BVALID),
    .m_axi_RDATA(m_axi_in_11_RDATA),
    .m_axi_RID(m_axi_in_11_RID),
    .m_axi_RLAST(m_axi_in_11_RLAST),
    .m_axi_RREADY(m_axi_in_11_RREADY),
    .m_axi_RRESP(m_axi_in_11_RRESP),
    .m_axi_RVALID(m_axi_in_11_RVALID),
    .m_axi_WDATA(m_axi_in_11_WDATA),
    .m_axi_WLAST(m_axi_in_11_WLAST),
    .m_axi_WREADY(m_axi_in_11_WREADY),
    .m_axi_WSTRB(m_axi_in_11_WSTRB),
    .m_axi_WVALID(m_axi_in_11_WVALID),
    .read_addr_din(in_11_read_addr__din),
    .read_addr_full_n(in_11_read_addr__full_n),
    .read_addr_write(in_11_read_addr__write),
    .read_data_dout(in_11_read_data__dout),
    .read_data_empty_n(in_11_read_data__empty_n),
    .read_data_read(in_11_read_data__read),
    .write_addr_din(in_11_write_addr__din),
    .write_addr_full_n(in_11_write_addr__full_n),
    .write_addr_write(in_11_write_addr__write),
    .write_data_din(in_11_write_data__din),
    .write_data_full_n(in_11_write_data__full_n),
    .write_data_write(in_11_write_data__write),
    .write_resp_dout(in_11_write_resp__dout),
    .write_resp_empty_n(in_11_write_resp__empty_n),
    .write_resp_read(in_11_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_11__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_11___out_11__q0),
    .m_axi_ARADDR(m_axi_out_11_ARADDR),
    .m_axi_ARBURST(m_axi_out_11_ARBURST),
    .m_axi_ARCACHE(m_axi_out_11_ARCACHE),
    .m_axi_ARID(m_axi_out_11_ARID),
    .m_axi_ARLEN(m_axi_out_11_ARLEN),
    .m_axi_ARLOCK(m_axi_out_11_ARLOCK),
    .m_axi_ARPROT(m_axi_out_11_ARPROT),
    .m_axi_ARQOS(m_axi_out_11_ARQOS),
    .m_axi_ARREADY(m_axi_out_11_ARREADY),
    .m_axi_ARSIZE(m_axi_out_11_ARSIZE),
    .m_axi_ARVALID(m_axi_out_11_ARVALID),
    .m_axi_AWADDR(m_axi_out_11_AWADDR),
    .m_axi_AWBURST(m_axi_out_11_AWBURST),
    .m_axi_AWCACHE(m_axi_out_11_AWCACHE),
    .m_axi_AWID(m_axi_out_11_AWID),
    .m_axi_AWLEN(m_axi_out_11_AWLEN),
    .m_axi_AWLOCK(m_axi_out_11_AWLOCK),
    .m_axi_AWPROT(m_axi_out_11_AWPROT),
    .m_axi_AWQOS(m_axi_out_11_AWQOS),
    .m_axi_AWREADY(m_axi_out_11_AWREADY),
    .m_axi_AWSIZE(m_axi_out_11_AWSIZE),
    .m_axi_AWVALID(m_axi_out_11_AWVALID),
    .m_axi_BID(m_axi_out_11_BID),
    .m_axi_BREADY(m_axi_out_11_BREADY),
    .m_axi_BRESP(m_axi_out_11_BRESP),
    .m_axi_BVALID(m_axi_out_11_BVALID),
    .m_axi_RDATA(m_axi_out_11_RDATA),
    .m_axi_RID(m_axi_out_11_RID),
    .m_axi_RLAST(m_axi_out_11_RLAST),
    .m_axi_RREADY(m_axi_out_11_RREADY),
    .m_axi_RRESP(m_axi_out_11_RRESP),
    .m_axi_RVALID(m_axi_out_11_RVALID),
    .m_axi_WDATA(m_axi_out_11_WDATA),
    .m_axi_WLAST(m_axi_out_11_WLAST),
    .m_axi_WREADY(m_axi_out_11_WREADY),
    .m_axi_WSTRB(m_axi_out_11_WSTRB),
    .m_axi_WVALID(m_axi_out_11_WVALID),
    .read_addr_din(out_11_read_addr__din),
    .read_addr_full_n(out_11_read_addr__full_n),
    .read_addr_write(out_11_read_addr__write),
    .read_data_dout(out_11_read_data__dout),
    .read_data_empty_n(out_11_read_data__empty_n),
    .read_data_read(out_11_read_data__read),
    .write_addr_din(out_11_write_addr__din),
    .write_addr_full_n(out_11_write_addr__full_n),
    .write_addr_write(out_11_write_addr__write),
    .write_data_din(out_11_write_data__din),
    .write_data_full_n(out_11_write_data__full_n),
    .write_data_write(out_11_write_data__write),
    .write_resp_dout(out_11_write_resp__dout),
    .write_resp_empty_n(out_11_write_resp__empty_n),
    .write_resp_read(out_11_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_12__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_12___in_12__q0),
    .m_axi_ARADDR(m_axi_in_12_ARADDR),
    .m_axi_ARBURST(m_axi_in_12_ARBURST),
    .m_axi_ARCACHE(m_axi_in_12_ARCACHE),
    .m_axi_ARID(m_axi_in_12_ARID),
    .m_axi_ARLEN(m_axi_in_12_ARLEN),
    .m_axi_ARLOCK(m_axi_in_12_ARLOCK),
    .m_axi_ARPROT(m_axi_in_12_ARPROT),
    .m_axi_ARQOS(m_axi_in_12_ARQOS),
    .m_axi_ARREADY(m_axi_in_12_ARREADY),
    .m_axi_ARSIZE(m_axi_in_12_ARSIZE),
    .m_axi_ARVALID(m_axi_in_12_ARVALID),
    .m_axi_AWADDR(m_axi_in_12_AWADDR),
    .m_axi_AWBURST(m_axi_in_12_AWBURST),
    .m_axi_AWCACHE(m_axi_in_12_AWCACHE),
    .m_axi_AWID(m_axi_in_12_AWID),
    .m_axi_AWLEN(m_axi_in_12_AWLEN),
    .m_axi_AWLOCK(m_axi_in_12_AWLOCK),
    .m_axi_AWPROT(m_axi_in_12_AWPROT),
    .m_axi_AWQOS(m_axi_in_12_AWQOS),
    .m_axi_AWREADY(m_axi_in_12_AWREADY),
    .m_axi_AWSIZE(m_axi_in_12_AWSIZE),
    .m_axi_AWVALID(m_axi_in_12_AWVALID),
    .m_axi_BID(m_axi_in_12_BID),
    .m_axi_BREADY(m_axi_in_12_BREADY),
    .m_axi_BRESP(m_axi_in_12_BRESP),
    .m_axi_BVALID(m_axi_in_12_BVALID),
    .m_axi_RDATA(m_axi_in_12_RDATA),
    .m_axi_RID(m_axi_in_12_RID),
    .m_axi_RLAST(m_axi_in_12_RLAST),
    .m_axi_RREADY(m_axi_in_12_RREADY),
    .m_axi_RRESP(m_axi_in_12_RRESP),
    .m_axi_RVALID(m_axi_in_12_RVALID),
    .m_axi_WDATA(m_axi_in_12_WDATA),
    .m_axi_WLAST(m_axi_in_12_WLAST),
    .m_axi_WREADY(m_axi_in_12_WREADY),
    .m_axi_WSTRB(m_axi_in_12_WSTRB),
    .m_axi_WVALID(m_axi_in_12_WVALID),
    .read_addr_din(in_12_read_addr__din),
    .read_addr_full_n(in_12_read_addr__full_n),
    .read_addr_write(in_12_read_addr__write),
    .read_data_dout(in_12_read_data__dout),
    .read_data_empty_n(in_12_read_data__empty_n),
    .read_data_read(in_12_read_data__read),
    .write_addr_din(in_12_write_addr__din),
    .write_addr_full_n(in_12_write_addr__full_n),
    .write_addr_write(in_12_write_addr__write),
    .write_data_din(in_12_write_data__din),
    .write_data_full_n(in_12_write_data__full_n),
    .write_data_write(in_12_write_data__write),
    .write_resp_dout(in_12_write_resp__dout),
    .write_resp_empty_n(in_12_write_resp__empty_n),
    .write_resp_read(in_12_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_12__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_12___out_12__q0),
    .m_axi_ARADDR(m_axi_out_12_ARADDR),
    .m_axi_ARBURST(m_axi_out_12_ARBURST),
    .m_axi_ARCACHE(m_axi_out_12_ARCACHE),
    .m_axi_ARID(m_axi_out_12_ARID),
    .m_axi_ARLEN(m_axi_out_12_ARLEN),
    .m_axi_ARLOCK(m_axi_out_12_ARLOCK),
    .m_axi_ARPROT(m_axi_out_12_ARPROT),
    .m_axi_ARQOS(m_axi_out_12_ARQOS),
    .m_axi_ARREADY(m_axi_out_12_ARREADY),
    .m_axi_ARSIZE(m_axi_out_12_ARSIZE),
    .m_axi_ARVALID(m_axi_out_12_ARVALID),
    .m_axi_AWADDR(m_axi_out_12_AWADDR),
    .m_axi_AWBURST(m_axi_out_12_AWBURST),
    .m_axi_AWCACHE(m_axi_out_12_AWCACHE),
    .m_axi_AWID(m_axi_out_12_AWID),
    .m_axi_AWLEN(m_axi_out_12_AWLEN),
    .m_axi_AWLOCK(m_axi_out_12_AWLOCK),
    .m_axi_AWPROT(m_axi_out_12_AWPROT),
    .m_axi_AWQOS(m_axi_out_12_AWQOS),
    .m_axi_AWREADY(m_axi_out_12_AWREADY),
    .m_axi_AWSIZE(m_axi_out_12_AWSIZE),
    .m_axi_AWVALID(m_axi_out_12_AWVALID),
    .m_axi_BID(m_axi_out_12_BID),
    .m_axi_BREADY(m_axi_out_12_BREADY),
    .m_axi_BRESP(m_axi_out_12_BRESP),
    .m_axi_BVALID(m_axi_out_12_BVALID),
    .m_axi_RDATA(m_axi_out_12_RDATA),
    .m_axi_RID(m_axi_out_12_RID),
    .m_axi_RLAST(m_axi_out_12_RLAST),
    .m_axi_RREADY(m_axi_out_12_RREADY),
    .m_axi_RRESP(m_axi_out_12_RRESP),
    .m_axi_RVALID(m_axi_out_12_RVALID),
    .m_axi_WDATA(m_axi_out_12_WDATA),
    .m_axi_WLAST(m_axi_out_12_WLAST),
    .m_axi_WREADY(m_axi_out_12_WREADY),
    .m_axi_WSTRB(m_axi_out_12_WSTRB),
    .m_axi_WVALID(m_axi_out_12_WVALID),
    .read_addr_din(out_12_read_addr__din),
    .read_addr_full_n(out_12_read_addr__full_n),
    .read_addr_write(out_12_read_addr__write),
    .read_data_dout(out_12_read_data__dout),
    .read_data_empty_n(out_12_read_data__empty_n),
    .read_data_read(out_12_read_data__read),
    .write_addr_din(out_12_write_addr__din),
    .write_addr_full_n(out_12_write_addr__full_n),
    .write_addr_write(out_12_write_addr__write),
    .write_data_din(out_12_write_data__din),
    .write_data_full_n(out_12_write_data__full_n),
    .write_data_write(out_12_write_data__write),
    .write_resp_dout(out_12_write_resp__dout),
    .write_resp_empty_n(out_12_write_resp__empty_n),
    .write_resp_read(out_12_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_13__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_13___in_13__q0),
    .m_axi_ARADDR(m_axi_in_13_ARADDR),
    .m_axi_ARBURST(m_axi_in_13_ARBURST),
    .m_axi_ARCACHE(m_axi_in_13_ARCACHE),
    .m_axi_ARID(m_axi_in_13_ARID),
    .m_axi_ARLEN(m_axi_in_13_ARLEN),
    .m_axi_ARLOCK(m_axi_in_13_ARLOCK),
    .m_axi_ARPROT(m_axi_in_13_ARPROT),
    .m_axi_ARQOS(m_axi_in_13_ARQOS),
    .m_axi_ARREADY(m_axi_in_13_ARREADY),
    .m_axi_ARSIZE(m_axi_in_13_ARSIZE),
    .m_axi_ARVALID(m_axi_in_13_ARVALID),
    .m_axi_AWADDR(m_axi_in_13_AWADDR),
    .m_axi_AWBURST(m_axi_in_13_AWBURST),
    .m_axi_AWCACHE(m_axi_in_13_AWCACHE),
    .m_axi_AWID(m_axi_in_13_AWID),
    .m_axi_AWLEN(m_axi_in_13_AWLEN),
    .m_axi_AWLOCK(m_axi_in_13_AWLOCK),
    .m_axi_AWPROT(m_axi_in_13_AWPROT),
    .m_axi_AWQOS(m_axi_in_13_AWQOS),
    .m_axi_AWREADY(m_axi_in_13_AWREADY),
    .m_axi_AWSIZE(m_axi_in_13_AWSIZE),
    .m_axi_AWVALID(m_axi_in_13_AWVALID),
    .m_axi_BID(m_axi_in_13_BID),
    .m_axi_BREADY(m_axi_in_13_BREADY),
    .m_axi_BRESP(m_axi_in_13_BRESP),
    .m_axi_BVALID(m_axi_in_13_BVALID),
    .m_axi_RDATA(m_axi_in_13_RDATA),
    .m_axi_RID(m_axi_in_13_RID),
    .m_axi_RLAST(m_axi_in_13_RLAST),
    .m_axi_RREADY(m_axi_in_13_RREADY),
    .m_axi_RRESP(m_axi_in_13_RRESP),
    .m_axi_RVALID(m_axi_in_13_RVALID),
    .m_axi_WDATA(m_axi_in_13_WDATA),
    .m_axi_WLAST(m_axi_in_13_WLAST),
    .m_axi_WREADY(m_axi_in_13_WREADY),
    .m_axi_WSTRB(m_axi_in_13_WSTRB),
    .m_axi_WVALID(m_axi_in_13_WVALID),
    .read_addr_din(in_13_read_addr__din),
    .read_addr_full_n(in_13_read_addr__full_n),
    .read_addr_write(in_13_read_addr__write),
    .read_data_dout(in_13_read_data__dout),
    .read_data_empty_n(in_13_read_data__empty_n),
    .read_data_read(in_13_read_data__read),
    .write_addr_din(in_13_write_addr__din),
    .write_addr_full_n(in_13_write_addr__full_n),
    .write_addr_write(in_13_write_addr__write),
    .write_data_din(in_13_write_data__din),
    .write_data_full_n(in_13_write_data__full_n),
    .write_data_write(in_13_write_data__write),
    .write_resp_dout(in_13_write_resp__dout),
    .write_resp_empty_n(in_13_write_resp__empty_n),
    .write_resp_read(in_13_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_13__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_13___out_13__q0),
    .m_axi_ARADDR(m_axi_out_13_ARADDR),
    .m_axi_ARBURST(m_axi_out_13_ARBURST),
    .m_axi_ARCACHE(m_axi_out_13_ARCACHE),
    .m_axi_ARID(m_axi_out_13_ARID),
    .m_axi_ARLEN(m_axi_out_13_ARLEN),
    .m_axi_ARLOCK(m_axi_out_13_ARLOCK),
    .m_axi_ARPROT(m_axi_out_13_ARPROT),
    .m_axi_ARQOS(m_axi_out_13_ARQOS),
    .m_axi_ARREADY(m_axi_out_13_ARREADY),
    .m_axi_ARSIZE(m_axi_out_13_ARSIZE),
    .m_axi_ARVALID(m_axi_out_13_ARVALID),
    .m_axi_AWADDR(m_axi_out_13_AWADDR),
    .m_axi_AWBURST(m_axi_out_13_AWBURST),
    .m_axi_AWCACHE(m_axi_out_13_AWCACHE),
    .m_axi_AWID(m_axi_out_13_AWID),
    .m_axi_AWLEN(m_axi_out_13_AWLEN),
    .m_axi_AWLOCK(m_axi_out_13_AWLOCK),
    .m_axi_AWPROT(m_axi_out_13_AWPROT),
    .m_axi_AWQOS(m_axi_out_13_AWQOS),
    .m_axi_AWREADY(m_axi_out_13_AWREADY),
    .m_axi_AWSIZE(m_axi_out_13_AWSIZE),
    .m_axi_AWVALID(m_axi_out_13_AWVALID),
    .m_axi_BID(m_axi_out_13_BID),
    .m_axi_BREADY(m_axi_out_13_BREADY),
    .m_axi_BRESP(m_axi_out_13_BRESP),
    .m_axi_BVALID(m_axi_out_13_BVALID),
    .m_axi_RDATA(m_axi_out_13_RDATA),
    .m_axi_RID(m_axi_out_13_RID),
    .m_axi_RLAST(m_axi_out_13_RLAST),
    .m_axi_RREADY(m_axi_out_13_RREADY),
    .m_axi_RRESP(m_axi_out_13_RRESP),
    .m_axi_RVALID(m_axi_out_13_RVALID),
    .m_axi_WDATA(m_axi_out_13_WDATA),
    .m_axi_WLAST(m_axi_out_13_WLAST),
    .m_axi_WREADY(m_axi_out_13_WREADY),
    .m_axi_WSTRB(m_axi_out_13_WSTRB),
    .m_axi_WVALID(m_axi_out_13_WVALID),
    .read_addr_din(out_13_read_addr__din),
    .read_addr_full_n(out_13_read_addr__full_n),
    .read_addr_write(out_13_read_addr__write),
    .read_data_dout(out_13_read_data__dout),
    .read_data_empty_n(out_13_read_data__empty_n),
    .read_data_read(out_13_read_data__read),
    .write_addr_din(out_13_write_addr__din),
    .write_addr_full_n(out_13_write_addr__full_n),
    .write_addr_write(out_13_write_addr__write),
    .write_data_din(out_13_write_data__din),
    .write_data_full_n(out_13_write_data__full_n),
    .write_data_write(out_13_write_data__write),
    .write_resp_dout(out_13_write_resp__dout),
    .write_resp_empty_n(out_13_write_resp__empty_n),
    .write_resp_read(out_13_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  in_14__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_14___in_14__q0),
    .m_axi_ARADDR(m_axi_in_14_ARADDR),
    .m_axi_ARBURST(m_axi_in_14_ARBURST),
    .m_axi_ARCACHE(m_axi_in_14_ARCACHE),
    .m_axi_ARID(m_axi_in_14_ARID),
    .m_axi_ARLEN(m_axi_in_14_ARLEN),
    .m_axi_ARLOCK(m_axi_in_14_ARLOCK),
    .m_axi_ARPROT(m_axi_in_14_ARPROT),
    .m_axi_ARQOS(m_axi_in_14_ARQOS),
    .m_axi_ARREADY(m_axi_in_14_ARREADY),
    .m_axi_ARSIZE(m_axi_in_14_ARSIZE),
    .m_axi_ARVALID(m_axi_in_14_ARVALID),
    .m_axi_AWADDR(m_axi_in_14_AWADDR),
    .m_axi_AWBURST(m_axi_in_14_AWBURST),
    .m_axi_AWCACHE(m_axi_in_14_AWCACHE),
    .m_axi_AWID(m_axi_in_14_AWID),
    .m_axi_AWLEN(m_axi_in_14_AWLEN),
    .m_axi_AWLOCK(m_axi_in_14_AWLOCK),
    .m_axi_AWPROT(m_axi_in_14_AWPROT),
    .m_axi_AWQOS(m_axi_in_14_AWQOS),
    .m_axi_AWREADY(m_axi_in_14_AWREADY),
    .m_axi_AWSIZE(m_axi_in_14_AWSIZE),
    .m_axi_AWVALID(m_axi_in_14_AWVALID),
    .m_axi_BID(m_axi_in_14_BID),
    .m_axi_BREADY(m_axi_in_14_BREADY),
    .m_axi_BRESP(m_axi_in_14_BRESP),
    .m_axi_BVALID(m_axi_in_14_BVALID),
    .m_axi_RDATA(m_axi_in_14_RDATA),
    .m_axi_RID(m_axi_in_14_RID),
    .m_axi_RLAST(m_axi_in_14_RLAST),
    .m_axi_RREADY(m_axi_in_14_RREADY),
    .m_axi_RRESP(m_axi_in_14_RRESP),
    .m_axi_RVALID(m_axi_in_14_RVALID),
    .m_axi_WDATA(m_axi_in_14_WDATA),
    .m_axi_WLAST(m_axi_in_14_WLAST),
    .m_axi_WREADY(m_axi_in_14_WREADY),
    .m_axi_WSTRB(m_axi_in_14_WSTRB),
    .m_axi_WVALID(m_axi_in_14_WVALID),
    .read_addr_din(in_14_read_addr__din),
    .read_addr_full_n(in_14_read_addr__full_n),
    .read_addr_write(in_14_read_addr__write),
    .read_data_dout(in_14_read_data__dout),
    .read_data_empty_n(in_14_read_data__empty_n),
    .read_data_read(in_14_read_data__read),
    .write_addr_din(in_14_write_addr__din),
    .write_addr_full_n(in_14_write_addr__full_n),
    .write_addr_write(in_14_write_addr__write),
    .write_data_din(in_14_write_data__din),
    .write_data_full_n(in_14_write_data__full_n),
    .write_data_write(in_14_write_data__write),
    .write_resp_dout(in_14_write_resp__dout),
    .write_resp_empty_n(in_14_write_resp__empty_n),
    .write_resp_read(in_14_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  out_14__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(inter_kernel_14___out_14__q0),
    .m_axi_ARADDR(m_axi_out_14_ARADDR),
    .m_axi_ARBURST(m_axi_out_14_ARBURST),
    .m_axi_ARCACHE(m_axi_out_14_ARCACHE),
    .m_axi_ARID(m_axi_out_14_ARID),
    .m_axi_ARLEN(m_axi_out_14_ARLEN),
    .m_axi_ARLOCK(m_axi_out_14_ARLOCK),
    .m_axi_ARPROT(m_axi_out_14_ARPROT),
    .m_axi_ARQOS(m_axi_out_14_ARQOS),
    .m_axi_ARREADY(m_axi_out_14_ARREADY),
    .m_axi_ARSIZE(m_axi_out_14_ARSIZE),
    .m_axi_ARVALID(m_axi_out_14_ARVALID),
    .m_axi_AWADDR(m_axi_out_14_AWADDR),
    .m_axi_AWBURST(m_axi_out_14_AWBURST),
    .m_axi_AWCACHE(m_axi_out_14_AWCACHE),
    .m_axi_AWID(m_axi_out_14_AWID),
    .m_axi_AWLEN(m_axi_out_14_AWLEN),
    .m_axi_AWLOCK(m_axi_out_14_AWLOCK),
    .m_axi_AWPROT(m_axi_out_14_AWPROT),
    .m_axi_AWQOS(m_axi_out_14_AWQOS),
    .m_axi_AWREADY(m_axi_out_14_AWREADY),
    .m_axi_AWSIZE(m_axi_out_14_AWSIZE),
    .m_axi_AWVALID(m_axi_out_14_AWVALID),
    .m_axi_BID(m_axi_out_14_BID),
    .m_axi_BREADY(m_axi_out_14_BREADY),
    .m_axi_BRESP(m_axi_out_14_BRESP),
    .m_axi_BVALID(m_axi_out_14_BVALID),
    .m_axi_RDATA(m_axi_out_14_RDATA),
    .m_axi_RID(m_axi_out_14_RID),
    .m_axi_RLAST(m_axi_out_14_RLAST),
    .m_axi_RREADY(m_axi_out_14_RREADY),
    .m_axi_RRESP(m_axi_out_14_RRESP),
    .m_axi_RVALID(m_axi_out_14_RVALID),
    .m_axi_WDATA(m_axi_out_14_WDATA),
    .m_axi_WLAST(m_axi_out_14_WLAST),
    .m_axi_WREADY(m_axi_out_14_WREADY),
    .m_axi_WSTRB(m_axi_out_14_WSTRB),
    .m_axi_WVALID(m_axi_out_14_WVALID),
    .read_addr_din(out_14_read_addr__din),
    .read_addr_full_n(out_14_read_addr__full_n),
    .read_addr_write(out_14_read_addr__write),
    .read_data_dout(out_14_read_data__dout),
    .read_data_empty_n(out_14_read_data__empty_n),
    .read_data_read(out_14_read_data__read),
    .write_addr_din(out_14_write_addr__din),
    .write_addr_full_n(out_14_write_addr__full_n),
    .write_addr_write(out_14_write_addr__write),
    .write_data_din(out_14_write_data__din),
    .write_data_full_n(out_14_write_data__full_n),
    .write_data_write(out_14_write_data__write),
    .write_resp_dout(out_14_write_resp__dout),
    .write_resp_empty_n(out_14_write_resp__empty_n),
    .write_resp_read(out_14_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) unikernel_fsm
  __tapa_fsm_unit
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .JACOBI3D_0__ap_start(JACOBI3D_0__ap_start),
    .JACOBI3D_0__ap_ready(JACOBI3D_0__ap_ready),
    .JACOBI3D_0__ap_done(JACOBI3D_0__ap_done),
    .JACOBI3D_0__ap_idle(JACOBI3D_0__ap_idle),
    .JACOBI3D_1__ap_start(JACOBI3D_1__ap_start),
    .JACOBI3D_1__ap_ready(JACOBI3D_1__ap_ready),
    .JACOBI3D_1__ap_done(JACOBI3D_1__ap_done),
    .JACOBI3D_1__ap_idle(JACOBI3D_1__ap_idle),
    .JACOBI3D_2__ap_start(JACOBI3D_2__ap_start),
    .JACOBI3D_2__ap_ready(JACOBI3D_2__ap_ready),
    .JACOBI3D_2__ap_done(JACOBI3D_2__ap_done),
    .JACOBI3D_2__ap_idle(JACOBI3D_2__ap_idle),
    .JACOBI3D_3__ap_start(JACOBI3D_3__ap_start),
    .JACOBI3D_3__ap_ready(JACOBI3D_3__ap_ready),
    .JACOBI3D_3__ap_done(JACOBI3D_3__ap_done),
    .JACOBI3D_3__ap_idle(JACOBI3D_3__ap_idle),
    .JACOBI3D_4__ap_start(JACOBI3D_4__ap_start),
    .JACOBI3D_4__ap_ready(JACOBI3D_4__ap_ready),
    .JACOBI3D_4__ap_done(JACOBI3D_4__ap_done),
    .JACOBI3D_4__ap_idle(JACOBI3D_4__ap_idle),
    .JACOBI3D_5__ap_start(JACOBI3D_5__ap_start),
    .JACOBI3D_5__ap_ready(JACOBI3D_5__ap_ready),
    .JACOBI3D_5__ap_done(JACOBI3D_5__ap_done),
    .JACOBI3D_5__ap_idle(JACOBI3D_5__ap_idle),
    .JACOBI3D_6__ap_start(JACOBI3D_6__ap_start),
    .JACOBI3D_6__ap_ready(JACOBI3D_6__ap_ready),
    .JACOBI3D_6__ap_done(JACOBI3D_6__ap_done),
    .JACOBI3D_6__ap_idle(JACOBI3D_6__ap_idle),
    .JACOBI3D_7__ap_start(JACOBI3D_7__ap_start),
    .JACOBI3D_7__ap_ready(JACOBI3D_7__ap_ready),
    .JACOBI3D_7__ap_done(JACOBI3D_7__ap_done),
    .JACOBI3D_7__ap_idle(JACOBI3D_7__ap_idle),
    .JACOBI3D_8__ap_start(JACOBI3D_8__ap_start),
    .JACOBI3D_8__ap_ready(JACOBI3D_8__ap_ready),
    .JACOBI3D_8__ap_done(JACOBI3D_8__ap_done),
    .JACOBI3D_8__ap_idle(JACOBI3D_8__ap_idle),
    .JACOBI3D_9__ap_start(JACOBI3D_9__ap_start),
    .JACOBI3D_9__ap_ready(JACOBI3D_9__ap_ready),
    .JACOBI3D_9__ap_done(JACOBI3D_9__ap_done),
    .JACOBI3D_9__ap_idle(JACOBI3D_9__ap_idle),
    .JACOBI3D_10__ap_start(JACOBI3D_10__ap_start),
    .JACOBI3D_10__ap_ready(JACOBI3D_10__ap_ready),
    .JACOBI3D_10__ap_done(JACOBI3D_10__ap_done),
    .JACOBI3D_10__ap_idle(JACOBI3D_10__ap_idle),
    .JACOBI3D_11__ap_start(JACOBI3D_11__ap_start),
    .JACOBI3D_11__ap_ready(JACOBI3D_11__ap_ready),
    .JACOBI3D_11__ap_done(JACOBI3D_11__ap_done),
    .JACOBI3D_11__ap_idle(JACOBI3D_11__ap_idle),
    .JACOBI3D_12__ap_start(JACOBI3D_12__ap_start),
    .JACOBI3D_12__ap_ready(JACOBI3D_12__ap_ready),
    .JACOBI3D_12__ap_done(JACOBI3D_12__ap_done),
    .JACOBI3D_12__ap_idle(JACOBI3D_12__ap_idle),
    .JACOBI3D_13__ap_start(JACOBI3D_13__ap_start),
    .JACOBI3D_13__ap_ready(JACOBI3D_13__ap_ready),
    .JACOBI3D_13__ap_done(JACOBI3D_13__ap_done),
    .JACOBI3D_13__ap_idle(JACOBI3D_13__ap_idle),
    .JACOBI3D_14__ap_start(JACOBI3D_14__ap_start),
    .JACOBI3D_14__ap_ready(JACOBI3D_14__ap_ready),
    .JACOBI3D_14__ap_done(JACOBI3D_14__ap_done),
    .JACOBI3D_14__ap_idle(JACOBI3D_14__ap_idle),
    .inter_kernel_0__ap_start(inter_kernel_0__ap_start),
    .inter_kernel_0__ap_ready(inter_kernel_0__ap_ready),
    .inter_kernel_0__ap_done(inter_kernel_0__ap_done),
    .inter_kernel_0__ap_idle(inter_kernel_0__ap_idle),
    .inter_kernel_1__ap_start(inter_kernel_1__ap_start),
    .inter_kernel_1__ap_ready(inter_kernel_1__ap_ready),
    .inter_kernel_1__ap_done(inter_kernel_1__ap_done),
    .inter_kernel_1__ap_idle(inter_kernel_1__ap_idle),
    .inter_kernel_2__ap_start(inter_kernel_2__ap_start),
    .inter_kernel_2__ap_ready(inter_kernel_2__ap_ready),
    .inter_kernel_2__ap_done(inter_kernel_2__ap_done),
    .inter_kernel_2__ap_idle(inter_kernel_2__ap_idle),
    .inter_kernel_3__ap_start(inter_kernel_3__ap_start),
    .inter_kernel_3__ap_ready(inter_kernel_3__ap_ready),
    .inter_kernel_3__ap_done(inter_kernel_3__ap_done),
    .inter_kernel_3__ap_idle(inter_kernel_3__ap_idle),
    .inter_kernel_4__ap_start(inter_kernel_4__ap_start),
    .inter_kernel_4__ap_ready(inter_kernel_4__ap_ready),
    .inter_kernel_4__ap_done(inter_kernel_4__ap_done),
    .inter_kernel_4__ap_idle(inter_kernel_4__ap_idle),
    .inter_kernel_5__ap_start(inter_kernel_5__ap_start),
    .inter_kernel_5__ap_ready(inter_kernel_5__ap_ready),
    .inter_kernel_5__ap_done(inter_kernel_5__ap_done),
    .inter_kernel_5__ap_idle(inter_kernel_5__ap_idle),
    .inter_kernel_6__ap_start(inter_kernel_6__ap_start),
    .inter_kernel_6__ap_ready(inter_kernel_6__ap_ready),
    .inter_kernel_6__ap_done(inter_kernel_6__ap_done),
    .inter_kernel_6__ap_idle(inter_kernel_6__ap_idle),
    .inter_kernel_7__ap_start(inter_kernel_7__ap_start),
    .inter_kernel_7__ap_ready(inter_kernel_7__ap_ready),
    .inter_kernel_7__ap_done(inter_kernel_7__ap_done),
    .inter_kernel_7__ap_idle(inter_kernel_7__ap_idle),
    .inter_kernel_8__ap_start(inter_kernel_8__ap_start),
    .inter_kernel_8__ap_ready(inter_kernel_8__ap_ready),
    .inter_kernel_8__ap_done(inter_kernel_8__ap_done),
    .inter_kernel_8__ap_idle(inter_kernel_8__ap_idle),
    .inter_kernel_9__ap_start(inter_kernel_9__ap_start),
    .inter_kernel_9__ap_ready(inter_kernel_9__ap_ready),
    .inter_kernel_9__ap_done(inter_kernel_9__ap_done),
    .inter_kernel_9__ap_idle(inter_kernel_9__ap_idle),
    .inter_kernel_10__ap_start(inter_kernel_10__ap_start),
    .inter_kernel_10__ap_ready(inter_kernel_10__ap_ready),
    .inter_kernel_10__ap_done(inter_kernel_10__ap_done),
    .inter_kernel_10__ap_idle(inter_kernel_10__ap_idle),
    .inter_kernel_11__ap_start(inter_kernel_11__ap_start),
    .inter_kernel_11__ap_ready(inter_kernel_11__ap_ready),
    .inter_kernel_11__ap_done(inter_kernel_11__ap_done),
    .inter_kernel_11__ap_idle(inter_kernel_11__ap_idle),
    .inter_kernel_12__ap_start(inter_kernel_12__ap_start),
    .inter_kernel_12__ap_ready(inter_kernel_12__ap_ready),
    .inter_kernel_12__ap_done(inter_kernel_12__ap_done),
    .inter_kernel_12__ap_idle(inter_kernel_12__ap_idle),
    .inter_kernel_13__ap_start(inter_kernel_13__ap_start),
    .inter_kernel_13__ap_ready(inter_kernel_13__ap_ready),
    .inter_kernel_13__ap_done(inter_kernel_13__ap_done),
    .inter_kernel_13__ap_idle(inter_kernel_13__ap_idle),
    .inter_kernel_14__ap_start(inter_kernel_14__ap_start),
    .inter_kernel_14__ap_ready(inter_kernel_14__ap_ready),
    .inter_kernel_14__ap_done(inter_kernel_14__ap_done),
    .inter_kernel_14__ap_idle(inter_kernel_14__ap_idle)
  );

  assign ap_rst_n_inv = (~ap_rst_n);
  assign JACOBI3D_0___iters__q0 = iters;
  assign JACOBI3D_1___iters__q0 = iters;
  assign JACOBI3D_2___iters__q0 = iters;
  assign JACOBI3D_3___iters__q0 = iters;
  assign JACOBI3D_4___iters__q0 = iters;
  assign JACOBI3D_5___iters__q0 = iters;
  assign JACOBI3D_6___iters__q0 = iters;
  assign JACOBI3D_7___iters__q0 = iters;
  assign JACOBI3D_8___iters__q0 = iters;
  assign JACOBI3D_9___iters__q0 = iters;
  assign JACOBI3D_10___iters__q0 = iters;
  assign JACOBI3D_11___iters__q0 = iters;
  assign JACOBI3D_12___iters__q0 = iters;
  assign JACOBI3D_13___iters__q0 = iters;
  assign JACOBI3D_14___iters__q0 = iters;
  assign inter_kernel_0___in_0__q0 = in_0;
  assign inter_kernel_0___iters__q0 = iters;
  assign inter_kernel_0___out_0__q0 = out_0;
  assign inter_kernel_1___in_1__q0 = in_1;
  assign inter_kernel_1___iters__q0 = iters;
  assign inter_kernel_1___out_1__q0 = out_1;
  assign inter_kernel_2___in_2__q0 = in_2;
  assign inter_kernel_2___iters__q0 = iters;
  assign inter_kernel_2___out_2__q0 = out_2;
  assign inter_kernel_3___in_3__q0 = in_3;
  assign inter_kernel_3___iters__q0 = iters;
  assign inter_kernel_3___out_3__q0 = out_3;
  assign inter_kernel_4___in_4__q0 = in_4;
  assign inter_kernel_4___iters__q0 = iters;
  assign inter_kernel_4___out_4__q0 = out_4;
  assign inter_kernel_5___in_5__q0 = in_5;
  assign inter_kernel_5___iters__q0 = iters;
  assign inter_kernel_5___out_5__q0 = out_5;
  assign inter_kernel_6___in_6__q0 = in_6;
  assign inter_kernel_6___iters__q0 = iters;
  assign inter_kernel_6___out_6__q0 = out_6;
  assign inter_kernel_7___in_7__q0 = in_7;
  assign inter_kernel_7___iters__q0 = iters;
  assign inter_kernel_7___out_7__q0 = out_7;
  assign inter_kernel_8___in_8__q0 = in_8;
  assign inter_kernel_8___iters__q0 = iters;
  assign inter_kernel_8___out_8__q0 = out_8;
  assign inter_kernel_9___in_9__q0 = in_9;
  assign inter_kernel_9___iters__q0 = iters;
  assign inter_kernel_9___out_9__q0 = out_9;
  assign inter_kernel_10___in_10__q0 = in_10;
  assign inter_kernel_10___iters__q0 = iters;
  assign inter_kernel_10___out_10__q0 = out_10;
  assign inter_kernel_11___in_11__q0 = in_11;
  assign inter_kernel_11___iters__q0 = iters;
  assign inter_kernel_11___out_11__q0 = out_11;
  assign inter_kernel_12___in_12__q0 = in_12;
  assign inter_kernel_12___iters__q0 = iters;
  assign inter_kernel_12___out_12__q0 = out_12;
  assign inter_kernel_13___in_13__q0 = in_13;
  assign inter_kernel_13___iters__q0 = iters;
  assign inter_kernel_13___out_13__q0 = out_13;
  assign inter_kernel_14___in_14__q0 = in_14;
  assign inter_kernel_14___iters__q0 = iters;
  assign inter_kernel_14___out_14__q0 = out_14;

endmodule
