`timescale 1 ns / 1 ps

(* CORE_GENERATION_INFO = "Sextans_Sextans,hls_ip_2022_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcu280-fsvh2892-2L-e,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2332,HLS_SYN_LUT=4200,HLS_VERSION=2022_2}" *)


module Sextans
(
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  ap_clk,
  ap_rst_n,
  interrupt,
  m_axi_edge_list_ch_0_ARADDR,
  m_axi_edge_list_ch_0_ARBURST,
  m_axi_edge_list_ch_0_ARCACHE,
  m_axi_edge_list_ch_0_ARID,
  m_axi_edge_list_ch_0_ARLEN,
  m_axi_edge_list_ch_0_ARLOCK,
  m_axi_edge_list_ch_0_ARPROT,
  m_axi_edge_list_ch_0_ARQOS,
  m_axi_edge_list_ch_0_ARREADY,
  m_axi_edge_list_ch_0_ARSIZE,
  m_axi_edge_list_ch_0_ARVALID,
  m_axi_edge_list_ch_0_AWADDR,
  m_axi_edge_list_ch_0_AWBURST,
  m_axi_edge_list_ch_0_AWCACHE,
  m_axi_edge_list_ch_0_AWID,
  m_axi_edge_list_ch_0_AWLEN,
  m_axi_edge_list_ch_0_AWLOCK,
  m_axi_edge_list_ch_0_AWPROT,
  m_axi_edge_list_ch_0_AWQOS,
  m_axi_edge_list_ch_0_AWREADY,
  m_axi_edge_list_ch_0_AWSIZE,
  m_axi_edge_list_ch_0_AWVALID,
  m_axi_edge_list_ch_0_BID,
  m_axi_edge_list_ch_0_BREADY,
  m_axi_edge_list_ch_0_BRESP,
  m_axi_edge_list_ch_0_BVALID,
  m_axi_edge_list_ch_0_RDATA,
  m_axi_edge_list_ch_0_RID,
  m_axi_edge_list_ch_0_RLAST,
  m_axi_edge_list_ch_0_RREADY,
  m_axi_edge_list_ch_0_RRESP,
  m_axi_edge_list_ch_0_RVALID,
  m_axi_edge_list_ch_0_WDATA,
  m_axi_edge_list_ch_0_WLAST,
  m_axi_edge_list_ch_0_WREADY,
  m_axi_edge_list_ch_0_WSTRB,
  m_axi_edge_list_ch_0_WVALID,
  m_axi_edge_list_ch_1_ARADDR,
  m_axi_edge_list_ch_1_ARBURST,
  m_axi_edge_list_ch_1_ARCACHE,
  m_axi_edge_list_ch_1_ARID,
  m_axi_edge_list_ch_1_ARLEN,
  m_axi_edge_list_ch_1_ARLOCK,
  m_axi_edge_list_ch_1_ARPROT,
  m_axi_edge_list_ch_1_ARQOS,
  m_axi_edge_list_ch_1_ARREADY,
  m_axi_edge_list_ch_1_ARSIZE,
  m_axi_edge_list_ch_1_ARVALID,
  m_axi_edge_list_ch_1_AWADDR,
  m_axi_edge_list_ch_1_AWBURST,
  m_axi_edge_list_ch_1_AWCACHE,
  m_axi_edge_list_ch_1_AWID,
  m_axi_edge_list_ch_1_AWLEN,
  m_axi_edge_list_ch_1_AWLOCK,
  m_axi_edge_list_ch_1_AWPROT,
  m_axi_edge_list_ch_1_AWQOS,
  m_axi_edge_list_ch_1_AWREADY,
  m_axi_edge_list_ch_1_AWSIZE,
  m_axi_edge_list_ch_1_AWVALID,
  m_axi_edge_list_ch_1_BID,
  m_axi_edge_list_ch_1_BREADY,
  m_axi_edge_list_ch_1_BRESP,
  m_axi_edge_list_ch_1_BVALID,
  m_axi_edge_list_ch_1_RDATA,
  m_axi_edge_list_ch_1_RID,
  m_axi_edge_list_ch_1_RLAST,
  m_axi_edge_list_ch_1_RREADY,
  m_axi_edge_list_ch_1_RRESP,
  m_axi_edge_list_ch_1_RVALID,
  m_axi_edge_list_ch_1_WDATA,
  m_axi_edge_list_ch_1_WLAST,
  m_axi_edge_list_ch_1_WREADY,
  m_axi_edge_list_ch_1_WSTRB,
  m_axi_edge_list_ch_1_WVALID,
  m_axi_edge_list_ch_2_ARADDR,
  m_axi_edge_list_ch_2_ARBURST,
  m_axi_edge_list_ch_2_ARCACHE,
  m_axi_edge_list_ch_2_ARID,
  m_axi_edge_list_ch_2_ARLEN,
  m_axi_edge_list_ch_2_ARLOCK,
  m_axi_edge_list_ch_2_ARPROT,
  m_axi_edge_list_ch_2_ARQOS,
  m_axi_edge_list_ch_2_ARREADY,
  m_axi_edge_list_ch_2_ARSIZE,
  m_axi_edge_list_ch_2_ARVALID,
  m_axi_edge_list_ch_2_AWADDR,
  m_axi_edge_list_ch_2_AWBURST,
  m_axi_edge_list_ch_2_AWCACHE,
  m_axi_edge_list_ch_2_AWID,
  m_axi_edge_list_ch_2_AWLEN,
  m_axi_edge_list_ch_2_AWLOCK,
  m_axi_edge_list_ch_2_AWPROT,
  m_axi_edge_list_ch_2_AWQOS,
  m_axi_edge_list_ch_2_AWREADY,
  m_axi_edge_list_ch_2_AWSIZE,
  m_axi_edge_list_ch_2_AWVALID,
  m_axi_edge_list_ch_2_BID,
  m_axi_edge_list_ch_2_BREADY,
  m_axi_edge_list_ch_2_BRESP,
  m_axi_edge_list_ch_2_BVALID,
  m_axi_edge_list_ch_2_RDATA,
  m_axi_edge_list_ch_2_RID,
  m_axi_edge_list_ch_2_RLAST,
  m_axi_edge_list_ch_2_RREADY,
  m_axi_edge_list_ch_2_RRESP,
  m_axi_edge_list_ch_2_RVALID,
  m_axi_edge_list_ch_2_WDATA,
  m_axi_edge_list_ch_2_WLAST,
  m_axi_edge_list_ch_2_WREADY,
  m_axi_edge_list_ch_2_WSTRB,
  m_axi_edge_list_ch_2_WVALID,
  m_axi_edge_list_ch_3_ARADDR,
  m_axi_edge_list_ch_3_ARBURST,
  m_axi_edge_list_ch_3_ARCACHE,
  m_axi_edge_list_ch_3_ARID,
  m_axi_edge_list_ch_3_ARLEN,
  m_axi_edge_list_ch_3_ARLOCK,
  m_axi_edge_list_ch_3_ARPROT,
  m_axi_edge_list_ch_3_ARQOS,
  m_axi_edge_list_ch_3_ARREADY,
  m_axi_edge_list_ch_3_ARSIZE,
  m_axi_edge_list_ch_3_ARVALID,
  m_axi_edge_list_ch_3_AWADDR,
  m_axi_edge_list_ch_3_AWBURST,
  m_axi_edge_list_ch_3_AWCACHE,
  m_axi_edge_list_ch_3_AWID,
  m_axi_edge_list_ch_3_AWLEN,
  m_axi_edge_list_ch_3_AWLOCK,
  m_axi_edge_list_ch_3_AWPROT,
  m_axi_edge_list_ch_3_AWQOS,
  m_axi_edge_list_ch_3_AWREADY,
  m_axi_edge_list_ch_3_AWSIZE,
  m_axi_edge_list_ch_3_AWVALID,
  m_axi_edge_list_ch_3_BID,
  m_axi_edge_list_ch_3_BREADY,
  m_axi_edge_list_ch_3_BRESP,
  m_axi_edge_list_ch_3_BVALID,
  m_axi_edge_list_ch_3_RDATA,
  m_axi_edge_list_ch_3_RID,
  m_axi_edge_list_ch_3_RLAST,
  m_axi_edge_list_ch_3_RREADY,
  m_axi_edge_list_ch_3_RRESP,
  m_axi_edge_list_ch_3_RVALID,
  m_axi_edge_list_ch_3_WDATA,
  m_axi_edge_list_ch_3_WLAST,
  m_axi_edge_list_ch_3_WREADY,
  m_axi_edge_list_ch_3_WSTRB,
  m_axi_edge_list_ch_3_WVALID,
  m_axi_edge_list_ch_4_ARADDR,
  m_axi_edge_list_ch_4_ARBURST,
  m_axi_edge_list_ch_4_ARCACHE,
  m_axi_edge_list_ch_4_ARID,
  m_axi_edge_list_ch_4_ARLEN,
  m_axi_edge_list_ch_4_ARLOCK,
  m_axi_edge_list_ch_4_ARPROT,
  m_axi_edge_list_ch_4_ARQOS,
  m_axi_edge_list_ch_4_ARREADY,
  m_axi_edge_list_ch_4_ARSIZE,
  m_axi_edge_list_ch_4_ARVALID,
  m_axi_edge_list_ch_4_AWADDR,
  m_axi_edge_list_ch_4_AWBURST,
  m_axi_edge_list_ch_4_AWCACHE,
  m_axi_edge_list_ch_4_AWID,
  m_axi_edge_list_ch_4_AWLEN,
  m_axi_edge_list_ch_4_AWLOCK,
  m_axi_edge_list_ch_4_AWPROT,
  m_axi_edge_list_ch_4_AWQOS,
  m_axi_edge_list_ch_4_AWREADY,
  m_axi_edge_list_ch_4_AWSIZE,
  m_axi_edge_list_ch_4_AWVALID,
  m_axi_edge_list_ch_4_BID,
  m_axi_edge_list_ch_4_BREADY,
  m_axi_edge_list_ch_4_BRESP,
  m_axi_edge_list_ch_4_BVALID,
  m_axi_edge_list_ch_4_RDATA,
  m_axi_edge_list_ch_4_RID,
  m_axi_edge_list_ch_4_RLAST,
  m_axi_edge_list_ch_4_RREADY,
  m_axi_edge_list_ch_4_RRESP,
  m_axi_edge_list_ch_4_RVALID,
  m_axi_edge_list_ch_4_WDATA,
  m_axi_edge_list_ch_4_WLAST,
  m_axi_edge_list_ch_4_WREADY,
  m_axi_edge_list_ch_4_WSTRB,
  m_axi_edge_list_ch_4_WVALID,
  m_axi_edge_list_ch_5_ARADDR,
  m_axi_edge_list_ch_5_ARBURST,
  m_axi_edge_list_ch_5_ARCACHE,
  m_axi_edge_list_ch_5_ARID,
  m_axi_edge_list_ch_5_ARLEN,
  m_axi_edge_list_ch_5_ARLOCK,
  m_axi_edge_list_ch_5_ARPROT,
  m_axi_edge_list_ch_5_ARQOS,
  m_axi_edge_list_ch_5_ARREADY,
  m_axi_edge_list_ch_5_ARSIZE,
  m_axi_edge_list_ch_5_ARVALID,
  m_axi_edge_list_ch_5_AWADDR,
  m_axi_edge_list_ch_5_AWBURST,
  m_axi_edge_list_ch_5_AWCACHE,
  m_axi_edge_list_ch_5_AWID,
  m_axi_edge_list_ch_5_AWLEN,
  m_axi_edge_list_ch_5_AWLOCK,
  m_axi_edge_list_ch_5_AWPROT,
  m_axi_edge_list_ch_5_AWQOS,
  m_axi_edge_list_ch_5_AWREADY,
  m_axi_edge_list_ch_5_AWSIZE,
  m_axi_edge_list_ch_5_AWVALID,
  m_axi_edge_list_ch_5_BID,
  m_axi_edge_list_ch_5_BREADY,
  m_axi_edge_list_ch_5_BRESP,
  m_axi_edge_list_ch_5_BVALID,
  m_axi_edge_list_ch_5_RDATA,
  m_axi_edge_list_ch_5_RID,
  m_axi_edge_list_ch_5_RLAST,
  m_axi_edge_list_ch_5_RREADY,
  m_axi_edge_list_ch_5_RRESP,
  m_axi_edge_list_ch_5_RVALID,
  m_axi_edge_list_ch_5_WDATA,
  m_axi_edge_list_ch_5_WLAST,
  m_axi_edge_list_ch_5_WREADY,
  m_axi_edge_list_ch_5_WSTRB,
  m_axi_edge_list_ch_5_WVALID,
  m_axi_edge_list_ch_6_ARADDR,
  m_axi_edge_list_ch_6_ARBURST,
  m_axi_edge_list_ch_6_ARCACHE,
  m_axi_edge_list_ch_6_ARID,
  m_axi_edge_list_ch_6_ARLEN,
  m_axi_edge_list_ch_6_ARLOCK,
  m_axi_edge_list_ch_6_ARPROT,
  m_axi_edge_list_ch_6_ARQOS,
  m_axi_edge_list_ch_6_ARREADY,
  m_axi_edge_list_ch_6_ARSIZE,
  m_axi_edge_list_ch_6_ARVALID,
  m_axi_edge_list_ch_6_AWADDR,
  m_axi_edge_list_ch_6_AWBURST,
  m_axi_edge_list_ch_6_AWCACHE,
  m_axi_edge_list_ch_6_AWID,
  m_axi_edge_list_ch_6_AWLEN,
  m_axi_edge_list_ch_6_AWLOCK,
  m_axi_edge_list_ch_6_AWPROT,
  m_axi_edge_list_ch_6_AWQOS,
  m_axi_edge_list_ch_6_AWREADY,
  m_axi_edge_list_ch_6_AWSIZE,
  m_axi_edge_list_ch_6_AWVALID,
  m_axi_edge_list_ch_6_BID,
  m_axi_edge_list_ch_6_BREADY,
  m_axi_edge_list_ch_6_BRESP,
  m_axi_edge_list_ch_6_BVALID,
  m_axi_edge_list_ch_6_RDATA,
  m_axi_edge_list_ch_6_RID,
  m_axi_edge_list_ch_6_RLAST,
  m_axi_edge_list_ch_6_RREADY,
  m_axi_edge_list_ch_6_RRESP,
  m_axi_edge_list_ch_6_RVALID,
  m_axi_edge_list_ch_6_WDATA,
  m_axi_edge_list_ch_6_WLAST,
  m_axi_edge_list_ch_6_WREADY,
  m_axi_edge_list_ch_6_WSTRB,
  m_axi_edge_list_ch_6_WVALID,
  m_axi_edge_list_ch_7_ARADDR,
  m_axi_edge_list_ch_7_ARBURST,
  m_axi_edge_list_ch_7_ARCACHE,
  m_axi_edge_list_ch_7_ARID,
  m_axi_edge_list_ch_7_ARLEN,
  m_axi_edge_list_ch_7_ARLOCK,
  m_axi_edge_list_ch_7_ARPROT,
  m_axi_edge_list_ch_7_ARQOS,
  m_axi_edge_list_ch_7_ARREADY,
  m_axi_edge_list_ch_7_ARSIZE,
  m_axi_edge_list_ch_7_ARVALID,
  m_axi_edge_list_ch_7_AWADDR,
  m_axi_edge_list_ch_7_AWBURST,
  m_axi_edge_list_ch_7_AWCACHE,
  m_axi_edge_list_ch_7_AWID,
  m_axi_edge_list_ch_7_AWLEN,
  m_axi_edge_list_ch_7_AWLOCK,
  m_axi_edge_list_ch_7_AWPROT,
  m_axi_edge_list_ch_7_AWQOS,
  m_axi_edge_list_ch_7_AWREADY,
  m_axi_edge_list_ch_7_AWSIZE,
  m_axi_edge_list_ch_7_AWVALID,
  m_axi_edge_list_ch_7_BID,
  m_axi_edge_list_ch_7_BREADY,
  m_axi_edge_list_ch_7_BRESP,
  m_axi_edge_list_ch_7_BVALID,
  m_axi_edge_list_ch_7_RDATA,
  m_axi_edge_list_ch_7_RID,
  m_axi_edge_list_ch_7_RLAST,
  m_axi_edge_list_ch_7_RREADY,
  m_axi_edge_list_ch_7_RRESP,
  m_axi_edge_list_ch_7_RVALID,
  m_axi_edge_list_ch_7_WDATA,
  m_axi_edge_list_ch_7_WLAST,
  m_axi_edge_list_ch_7_WREADY,
  m_axi_edge_list_ch_7_WSTRB,
  m_axi_edge_list_ch_7_WVALID,
  m_axi_mat_B_ch_0_ARADDR,
  m_axi_mat_B_ch_0_ARBURST,
  m_axi_mat_B_ch_0_ARCACHE,
  m_axi_mat_B_ch_0_ARID,
  m_axi_mat_B_ch_0_ARLEN,
  m_axi_mat_B_ch_0_ARLOCK,
  m_axi_mat_B_ch_0_ARPROT,
  m_axi_mat_B_ch_0_ARQOS,
  m_axi_mat_B_ch_0_ARREADY,
  m_axi_mat_B_ch_0_ARSIZE,
  m_axi_mat_B_ch_0_ARVALID,
  m_axi_mat_B_ch_0_AWADDR,
  m_axi_mat_B_ch_0_AWBURST,
  m_axi_mat_B_ch_0_AWCACHE,
  m_axi_mat_B_ch_0_AWID,
  m_axi_mat_B_ch_0_AWLEN,
  m_axi_mat_B_ch_0_AWLOCK,
  m_axi_mat_B_ch_0_AWPROT,
  m_axi_mat_B_ch_0_AWQOS,
  m_axi_mat_B_ch_0_AWREADY,
  m_axi_mat_B_ch_0_AWSIZE,
  m_axi_mat_B_ch_0_AWVALID,
  m_axi_mat_B_ch_0_BID,
  m_axi_mat_B_ch_0_BREADY,
  m_axi_mat_B_ch_0_BRESP,
  m_axi_mat_B_ch_0_BVALID,
  m_axi_mat_B_ch_0_RDATA,
  m_axi_mat_B_ch_0_RID,
  m_axi_mat_B_ch_0_RLAST,
  m_axi_mat_B_ch_0_RREADY,
  m_axi_mat_B_ch_0_RRESP,
  m_axi_mat_B_ch_0_RVALID,
  m_axi_mat_B_ch_0_WDATA,
  m_axi_mat_B_ch_0_WLAST,
  m_axi_mat_B_ch_0_WREADY,
  m_axi_mat_B_ch_0_WSTRB,
  m_axi_mat_B_ch_0_WVALID,
  m_axi_mat_B_ch_1_ARADDR,
  m_axi_mat_B_ch_1_ARBURST,
  m_axi_mat_B_ch_1_ARCACHE,
  m_axi_mat_B_ch_1_ARID,
  m_axi_mat_B_ch_1_ARLEN,
  m_axi_mat_B_ch_1_ARLOCK,
  m_axi_mat_B_ch_1_ARPROT,
  m_axi_mat_B_ch_1_ARQOS,
  m_axi_mat_B_ch_1_ARREADY,
  m_axi_mat_B_ch_1_ARSIZE,
  m_axi_mat_B_ch_1_ARVALID,
  m_axi_mat_B_ch_1_AWADDR,
  m_axi_mat_B_ch_1_AWBURST,
  m_axi_mat_B_ch_1_AWCACHE,
  m_axi_mat_B_ch_1_AWID,
  m_axi_mat_B_ch_1_AWLEN,
  m_axi_mat_B_ch_1_AWLOCK,
  m_axi_mat_B_ch_1_AWPROT,
  m_axi_mat_B_ch_1_AWQOS,
  m_axi_mat_B_ch_1_AWREADY,
  m_axi_mat_B_ch_1_AWSIZE,
  m_axi_mat_B_ch_1_AWVALID,
  m_axi_mat_B_ch_1_BID,
  m_axi_mat_B_ch_1_BREADY,
  m_axi_mat_B_ch_1_BRESP,
  m_axi_mat_B_ch_1_BVALID,
  m_axi_mat_B_ch_1_RDATA,
  m_axi_mat_B_ch_1_RID,
  m_axi_mat_B_ch_1_RLAST,
  m_axi_mat_B_ch_1_RREADY,
  m_axi_mat_B_ch_1_RRESP,
  m_axi_mat_B_ch_1_RVALID,
  m_axi_mat_B_ch_1_WDATA,
  m_axi_mat_B_ch_1_WLAST,
  m_axi_mat_B_ch_1_WREADY,
  m_axi_mat_B_ch_1_WSTRB,
  m_axi_mat_B_ch_1_WVALID,
  m_axi_mat_B_ch_2_ARADDR,
  m_axi_mat_B_ch_2_ARBURST,
  m_axi_mat_B_ch_2_ARCACHE,
  m_axi_mat_B_ch_2_ARID,
  m_axi_mat_B_ch_2_ARLEN,
  m_axi_mat_B_ch_2_ARLOCK,
  m_axi_mat_B_ch_2_ARPROT,
  m_axi_mat_B_ch_2_ARQOS,
  m_axi_mat_B_ch_2_ARREADY,
  m_axi_mat_B_ch_2_ARSIZE,
  m_axi_mat_B_ch_2_ARVALID,
  m_axi_mat_B_ch_2_AWADDR,
  m_axi_mat_B_ch_2_AWBURST,
  m_axi_mat_B_ch_2_AWCACHE,
  m_axi_mat_B_ch_2_AWID,
  m_axi_mat_B_ch_2_AWLEN,
  m_axi_mat_B_ch_2_AWLOCK,
  m_axi_mat_B_ch_2_AWPROT,
  m_axi_mat_B_ch_2_AWQOS,
  m_axi_mat_B_ch_2_AWREADY,
  m_axi_mat_B_ch_2_AWSIZE,
  m_axi_mat_B_ch_2_AWVALID,
  m_axi_mat_B_ch_2_BID,
  m_axi_mat_B_ch_2_BREADY,
  m_axi_mat_B_ch_2_BRESP,
  m_axi_mat_B_ch_2_BVALID,
  m_axi_mat_B_ch_2_RDATA,
  m_axi_mat_B_ch_2_RID,
  m_axi_mat_B_ch_2_RLAST,
  m_axi_mat_B_ch_2_RREADY,
  m_axi_mat_B_ch_2_RRESP,
  m_axi_mat_B_ch_2_RVALID,
  m_axi_mat_B_ch_2_WDATA,
  m_axi_mat_B_ch_2_WLAST,
  m_axi_mat_B_ch_2_WREADY,
  m_axi_mat_B_ch_2_WSTRB,
  m_axi_mat_B_ch_2_WVALID,
  m_axi_mat_B_ch_3_ARADDR,
  m_axi_mat_B_ch_3_ARBURST,
  m_axi_mat_B_ch_3_ARCACHE,
  m_axi_mat_B_ch_3_ARID,
  m_axi_mat_B_ch_3_ARLEN,
  m_axi_mat_B_ch_3_ARLOCK,
  m_axi_mat_B_ch_3_ARPROT,
  m_axi_mat_B_ch_3_ARQOS,
  m_axi_mat_B_ch_3_ARREADY,
  m_axi_mat_B_ch_3_ARSIZE,
  m_axi_mat_B_ch_3_ARVALID,
  m_axi_mat_B_ch_3_AWADDR,
  m_axi_mat_B_ch_3_AWBURST,
  m_axi_mat_B_ch_3_AWCACHE,
  m_axi_mat_B_ch_3_AWID,
  m_axi_mat_B_ch_3_AWLEN,
  m_axi_mat_B_ch_3_AWLOCK,
  m_axi_mat_B_ch_3_AWPROT,
  m_axi_mat_B_ch_3_AWQOS,
  m_axi_mat_B_ch_3_AWREADY,
  m_axi_mat_B_ch_3_AWSIZE,
  m_axi_mat_B_ch_3_AWVALID,
  m_axi_mat_B_ch_3_BID,
  m_axi_mat_B_ch_3_BREADY,
  m_axi_mat_B_ch_3_BRESP,
  m_axi_mat_B_ch_3_BVALID,
  m_axi_mat_B_ch_3_RDATA,
  m_axi_mat_B_ch_3_RID,
  m_axi_mat_B_ch_3_RLAST,
  m_axi_mat_B_ch_3_RREADY,
  m_axi_mat_B_ch_3_RRESP,
  m_axi_mat_B_ch_3_RVALID,
  m_axi_mat_B_ch_3_WDATA,
  m_axi_mat_B_ch_3_WLAST,
  m_axi_mat_B_ch_3_WREADY,
  m_axi_mat_B_ch_3_WSTRB,
  m_axi_mat_B_ch_3_WVALID,
  m_axi_mat_C_ch_in_0_ARADDR,
  m_axi_mat_C_ch_in_0_ARBURST,
  m_axi_mat_C_ch_in_0_ARCACHE,
  m_axi_mat_C_ch_in_0_ARID,
  m_axi_mat_C_ch_in_0_ARLEN,
  m_axi_mat_C_ch_in_0_ARLOCK,
  m_axi_mat_C_ch_in_0_ARPROT,
  m_axi_mat_C_ch_in_0_ARQOS,
  m_axi_mat_C_ch_in_0_ARREADY,
  m_axi_mat_C_ch_in_0_ARSIZE,
  m_axi_mat_C_ch_in_0_ARVALID,
  m_axi_mat_C_ch_in_0_AWADDR,
  m_axi_mat_C_ch_in_0_AWBURST,
  m_axi_mat_C_ch_in_0_AWCACHE,
  m_axi_mat_C_ch_in_0_AWID,
  m_axi_mat_C_ch_in_0_AWLEN,
  m_axi_mat_C_ch_in_0_AWLOCK,
  m_axi_mat_C_ch_in_0_AWPROT,
  m_axi_mat_C_ch_in_0_AWQOS,
  m_axi_mat_C_ch_in_0_AWREADY,
  m_axi_mat_C_ch_in_0_AWSIZE,
  m_axi_mat_C_ch_in_0_AWVALID,
  m_axi_mat_C_ch_in_0_BID,
  m_axi_mat_C_ch_in_0_BREADY,
  m_axi_mat_C_ch_in_0_BRESP,
  m_axi_mat_C_ch_in_0_BVALID,
  m_axi_mat_C_ch_in_0_RDATA,
  m_axi_mat_C_ch_in_0_RID,
  m_axi_mat_C_ch_in_0_RLAST,
  m_axi_mat_C_ch_in_0_RREADY,
  m_axi_mat_C_ch_in_0_RRESP,
  m_axi_mat_C_ch_in_0_RVALID,
  m_axi_mat_C_ch_in_0_WDATA,
  m_axi_mat_C_ch_in_0_WLAST,
  m_axi_mat_C_ch_in_0_WREADY,
  m_axi_mat_C_ch_in_0_WSTRB,
  m_axi_mat_C_ch_in_0_WVALID,
  m_axi_mat_C_ch_in_1_ARADDR,
  m_axi_mat_C_ch_in_1_ARBURST,
  m_axi_mat_C_ch_in_1_ARCACHE,
  m_axi_mat_C_ch_in_1_ARID,
  m_axi_mat_C_ch_in_1_ARLEN,
  m_axi_mat_C_ch_in_1_ARLOCK,
  m_axi_mat_C_ch_in_1_ARPROT,
  m_axi_mat_C_ch_in_1_ARQOS,
  m_axi_mat_C_ch_in_1_ARREADY,
  m_axi_mat_C_ch_in_1_ARSIZE,
  m_axi_mat_C_ch_in_1_ARVALID,
  m_axi_mat_C_ch_in_1_AWADDR,
  m_axi_mat_C_ch_in_1_AWBURST,
  m_axi_mat_C_ch_in_1_AWCACHE,
  m_axi_mat_C_ch_in_1_AWID,
  m_axi_mat_C_ch_in_1_AWLEN,
  m_axi_mat_C_ch_in_1_AWLOCK,
  m_axi_mat_C_ch_in_1_AWPROT,
  m_axi_mat_C_ch_in_1_AWQOS,
  m_axi_mat_C_ch_in_1_AWREADY,
  m_axi_mat_C_ch_in_1_AWSIZE,
  m_axi_mat_C_ch_in_1_AWVALID,
  m_axi_mat_C_ch_in_1_BID,
  m_axi_mat_C_ch_in_1_BREADY,
  m_axi_mat_C_ch_in_1_BRESP,
  m_axi_mat_C_ch_in_1_BVALID,
  m_axi_mat_C_ch_in_1_RDATA,
  m_axi_mat_C_ch_in_1_RID,
  m_axi_mat_C_ch_in_1_RLAST,
  m_axi_mat_C_ch_in_1_RREADY,
  m_axi_mat_C_ch_in_1_RRESP,
  m_axi_mat_C_ch_in_1_RVALID,
  m_axi_mat_C_ch_in_1_WDATA,
  m_axi_mat_C_ch_in_1_WLAST,
  m_axi_mat_C_ch_in_1_WREADY,
  m_axi_mat_C_ch_in_1_WSTRB,
  m_axi_mat_C_ch_in_1_WVALID,
  m_axi_mat_C_ch_in_2_ARADDR,
  m_axi_mat_C_ch_in_2_ARBURST,
  m_axi_mat_C_ch_in_2_ARCACHE,
  m_axi_mat_C_ch_in_2_ARID,
  m_axi_mat_C_ch_in_2_ARLEN,
  m_axi_mat_C_ch_in_2_ARLOCK,
  m_axi_mat_C_ch_in_2_ARPROT,
  m_axi_mat_C_ch_in_2_ARQOS,
  m_axi_mat_C_ch_in_2_ARREADY,
  m_axi_mat_C_ch_in_2_ARSIZE,
  m_axi_mat_C_ch_in_2_ARVALID,
  m_axi_mat_C_ch_in_2_AWADDR,
  m_axi_mat_C_ch_in_2_AWBURST,
  m_axi_mat_C_ch_in_2_AWCACHE,
  m_axi_mat_C_ch_in_2_AWID,
  m_axi_mat_C_ch_in_2_AWLEN,
  m_axi_mat_C_ch_in_2_AWLOCK,
  m_axi_mat_C_ch_in_2_AWPROT,
  m_axi_mat_C_ch_in_2_AWQOS,
  m_axi_mat_C_ch_in_2_AWREADY,
  m_axi_mat_C_ch_in_2_AWSIZE,
  m_axi_mat_C_ch_in_2_AWVALID,
  m_axi_mat_C_ch_in_2_BID,
  m_axi_mat_C_ch_in_2_BREADY,
  m_axi_mat_C_ch_in_2_BRESP,
  m_axi_mat_C_ch_in_2_BVALID,
  m_axi_mat_C_ch_in_2_RDATA,
  m_axi_mat_C_ch_in_2_RID,
  m_axi_mat_C_ch_in_2_RLAST,
  m_axi_mat_C_ch_in_2_RREADY,
  m_axi_mat_C_ch_in_2_RRESP,
  m_axi_mat_C_ch_in_2_RVALID,
  m_axi_mat_C_ch_in_2_WDATA,
  m_axi_mat_C_ch_in_2_WLAST,
  m_axi_mat_C_ch_in_2_WREADY,
  m_axi_mat_C_ch_in_2_WSTRB,
  m_axi_mat_C_ch_in_2_WVALID,
  m_axi_mat_C_ch_in_3_ARADDR,
  m_axi_mat_C_ch_in_3_ARBURST,
  m_axi_mat_C_ch_in_3_ARCACHE,
  m_axi_mat_C_ch_in_3_ARID,
  m_axi_mat_C_ch_in_3_ARLEN,
  m_axi_mat_C_ch_in_3_ARLOCK,
  m_axi_mat_C_ch_in_3_ARPROT,
  m_axi_mat_C_ch_in_3_ARQOS,
  m_axi_mat_C_ch_in_3_ARREADY,
  m_axi_mat_C_ch_in_3_ARSIZE,
  m_axi_mat_C_ch_in_3_ARVALID,
  m_axi_mat_C_ch_in_3_AWADDR,
  m_axi_mat_C_ch_in_3_AWBURST,
  m_axi_mat_C_ch_in_3_AWCACHE,
  m_axi_mat_C_ch_in_3_AWID,
  m_axi_mat_C_ch_in_3_AWLEN,
  m_axi_mat_C_ch_in_3_AWLOCK,
  m_axi_mat_C_ch_in_3_AWPROT,
  m_axi_mat_C_ch_in_3_AWQOS,
  m_axi_mat_C_ch_in_3_AWREADY,
  m_axi_mat_C_ch_in_3_AWSIZE,
  m_axi_mat_C_ch_in_3_AWVALID,
  m_axi_mat_C_ch_in_3_BID,
  m_axi_mat_C_ch_in_3_BREADY,
  m_axi_mat_C_ch_in_3_BRESP,
  m_axi_mat_C_ch_in_3_BVALID,
  m_axi_mat_C_ch_in_3_RDATA,
  m_axi_mat_C_ch_in_3_RID,
  m_axi_mat_C_ch_in_3_RLAST,
  m_axi_mat_C_ch_in_3_RREADY,
  m_axi_mat_C_ch_in_3_RRESP,
  m_axi_mat_C_ch_in_3_RVALID,
  m_axi_mat_C_ch_in_3_WDATA,
  m_axi_mat_C_ch_in_3_WLAST,
  m_axi_mat_C_ch_in_3_WREADY,
  m_axi_mat_C_ch_in_3_WSTRB,
  m_axi_mat_C_ch_in_3_WVALID,
  m_axi_mat_C_ch_in_4_ARADDR,
  m_axi_mat_C_ch_in_4_ARBURST,
  m_axi_mat_C_ch_in_4_ARCACHE,
  m_axi_mat_C_ch_in_4_ARID,
  m_axi_mat_C_ch_in_4_ARLEN,
  m_axi_mat_C_ch_in_4_ARLOCK,
  m_axi_mat_C_ch_in_4_ARPROT,
  m_axi_mat_C_ch_in_4_ARQOS,
  m_axi_mat_C_ch_in_4_ARREADY,
  m_axi_mat_C_ch_in_4_ARSIZE,
  m_axi_mat_C_ch_in_4_ARVALID,
  m_axi_mat_C_ch_in_4_AWADDR,
  m_axi_mat_C_ch_in_4_AWBURST,
  m_axi_mat_C_ch_in_4_AWCACHE,
  m_axi_mat_C_ch_in_4_AWID,
  m_axi_mat_C_ch_in_4_AWLEN,
  m_axi_mat_C_ch_in_4_AWLOCK,
  m_axi_mat_C_ch_in_4_AWPROT,
  m_axi_mat_C_ch_in_4_AWQOS,
  m_axi_mat_C_ch_in_4_AWREADY,
  m_axi_mat_C_ch_in_4_AWSIZE,
  m_axi_mat_C_ch_in_4_AWVALID,
  m_axi_mat_C_ch_in_4_BID,
  m_axi_mat_C_ch_in_4_BREADY,
  m_axi_mat_C_ch_in_4_BRESP,
  m_axi_mat_C_ch_in_4_BVALID,
  m_axi_mat_C_ch_in_4_RDATA,
  m_axi_mat_C_ch_in_4_RID,
  m_axi_mat_C_ch_in_4_RLAST,
  m_axi_mat_C_ch_in_4_RREADY,
  m_axi_mat_C_ch_in_4_RRESP,
  m_axi_mat_C_ch_in_4_RVALID,
  m_axi_mat_C_ch_in_4_WDATA,
  m_axi_mat_C_ch_in_4_WLAST,
  m_axi_mat_C_ch_in_4_WREADY,
  m_axi_mat_C_ch_in_4_WSTRB,
  m_axi_mat_C_ch_in_4_WVALID,
  m_axi_mat_C_ch_in_5_ARADDR,
  m_axi_mat_C_ch_in_5_ARBURST,
  m_axi_mat_C_ch_in_5_ARCACHE,
  m_axi_mat_C_ch_in_5_ARID,
  m_axi_mat_C_ch_in_5_ARLEN,
  m_axi_mat_C_ch_in_5_ARLOCK,
  m_axi_mat_C_ch_in_5_ARPROT,
  m_axi_mat_C_ch_in_5_ARQOS,
  m_axi_mat_C_ch_in_5_ARREADY,
  m_axi_mat_C_ch_in_5_ARSIZE,
  m_axi_mat_C_ch_in_5_ARVALID,
  m_axi_mat_C_ch_in_5_AWADDR,
  m_axi_mat_C_ch_in_5_AWBURST,
  m_axi_mat_C_ch_in_5_AWCACHE,
  m_axi_mat_C_ch_in_5_AWID,
  m_axi_mat_C_ch_in_5_AWLEN,
  m_axi_mat_C_ch_in_5_AWLOCK,
  m_axi_mat_C_ch_in_5_AWPROT,
  m_axi_mat_C_ch_in_5_AWQOS,
  m_axi_mat_C_ch_in_5_AWREADY,
  m_axi_mat_C_ch_in_5_AWSIZE,
  m_axi_mat_C_ch_in_5_AWVALID,
  m_axi_mat_C_ch_in_5_BID,
  m_axi_mat_C_ch_in_5_BREADY,
  m_axi_mat_C_ch_in_5_BRESP,
  m_axi_mat_C_ch_in_5_BVALID,
  m_axi_mat_C_ch_in_5_RDATA,
  m_axi_mat_C_ch_in_5_RID,
  m_axi_mat_C_ch_in_5_RLAST,
  m_axi_mat_C_ch_in_5_RREADY,
  m_axi_mat_C_ch_in_5_RRESP,
  m_axi_mat_C_ch_in_5_RVALID,
  m_axi_mat_C_ch_in_5_WDATA,
  m_axi_mat_C_ch_in_5_WLAST,
  m_axi_mat_C_ch_in_5_WREADY,
  m_axi_mat_C_ch_in_5_WSTRB,
  m_axi_mat_C_ch_in_5_WVALID,
  m_axi_mat_C_ch_in_6_ARADDR,
  m_axi_mat_C_ch_in_6_ARBURST,
  m_axi_mat_C_ch_in_6_ARCACHE,
  m_axi_mat_C_ch_in_6_ARID,
  m_axi_mat_C_ch_in_6_ARLEN,
  m_axi_mat_C_ch_in_6_ARLOCK,
  m_axi_mat_C_ch_in_6_ARPROT,
  m_axi_mat_C_ch_in_6_ARQOS,
  m_axi_mat_C_ch_in_6_ARREADY,
  m_axi_mat_C_ch_in_6_ARSIZE,
  m_axi_mat_C_ch_in_6_ARVALID,
  m_axi_mat_C_ch_in_6_AWADDR,
  m_axi_mat_C_ch_in_6_AWBURST,
  m_axi_mat_C_ch_in_6_AWCACHE,
  m_axi_mat_C_ch_in_6_AWID,
  m_axi_mat_C_ch_in_6_AWLEN,
  m_axi_mat_C_ch_in_6_AWLOCK,
  m_axi_mat_C_ch_in_6_AWPROT,
  m_axi_mat_C_ch_in_6_AWQOS,
  m_axi_mat_C_ch_in_6_AWREADY,
  m_axi_mat_C_ch_in_6_AWSIZE,
  m_axi_mat_C_ch_in_6_AWVALID,
  m_axi_mat_C_ch_in_6_BID,
  m_axi_mat_C_ch_in_6_BREADY,
  m_axi_mat_C_ch_in_6_BRESP,
  m_axi_mat_C_ch_in_6_BVALID,
  m_axi_mat_C_ch_in_6_RDATA,
  m_axi_mat_C_ch_in_6_RID,
  m_axi_mat_C_ch_in_6_RLAST,
  m_axi_mat_C_ch_in_6_RREADY,
  m_axi_mat_C_ch_in_6_RRESP,
  m_axi_mat_C_ch_in_6_RVALID,
  m_axi_mat_C_ch_in_6_WDATA,
  m_axi_mat_C_ch_in_6_WLAST,
  m_axi_mat_C_ch_in_6_WREADY,
  m_axi_mat_C_ch_in_6_WSTRB,
  m_axi_mat_C_ch_in_6_WVALID,
  m_axi_mat_C_ch_in_7_ARADDR,
  m_axi_mat_C_ch_in_7_ARBURST,
  m_axi_mat_C_ch_in_7_ARCACHE,
  m_axi_mat_C_ch_in_7_ARID,
  m_axi_mat_C_ch_in_7_ARLEN,
  m_axi_mat_C_ch_in_7_ARLOCK,
  m_axi_mat_C_ch_in_7_ARPROT,
  m_axi_mat_C_ch_in_7_ARQOS,
  m_axi_mat_C_ch_in_7_ARREADY,
  m_axi_mat_C_ch_in_7_ARSIZE,
  m_axi_mat_C_ch_in_7_ARVALID,
  m_axi_mat_C_ch_in_7_AWADDR,
  m_axi_mat_C_ch_in_7_AWBURST,
  m_axi_mat_C_ch_in_7_AWCACHE,
  m_axi_mat_C_ch_in_7_AWID,
  m_axi_mat_C_ch_in_7_AWLEN,
  m_axi_mat_C_ch_in_7_AWLOCK,
  m_axi_mat_C_ch_in_7_AWPROT,
  m_axi_mat_C_ch_in_7_AWQOS,
  m_axi_mat_C_ch_in_7_AWREADY,
  m_axi_mat_C_ch_in_7_AWSIZE,
  m_axi_mat_C_ch_in_7_AWVALID,
  m_axi_mat_C_ch_in_7_BID,
  m_axi_mat_C_ch_in_7_BREADY,
  m_axi_mat_C_ch_in_7_BRESP,
  m_axi_mat_C_ch_in_7_BVALID,
  m_axi_mat_C_ch_in_7_RDATA,
  m_axi_mat_C_ch_in_7_RID,
  m_axi_mat_C_ch_in_7_RLAST,
  m_axi_mat_C_ch_in_7_RREADY,
  m_axi_mat_C_ch_in_7_RRESP,
  m_axi_mat_C_ch_in_7_RVALID,
  m_axi_mat_C_ch_in_7_WDATA,
  m_axi_mat_C_ch_in_7_WLAST,
  m_axi_mat_C_ch_in_7_WREADY,
  m_axi_mat_C_ch_in_7_WSTRB,
  m_axi_mat_C_ch_in_7_WVALID,
  m_axi_edge_list_ptr_ARADDR,
  m_axi_edge_list_ptr_ARBURST,
  m_axi_edge_list_ptr_ARCACHE,
  m_axi_edge_list_ptr_ARID,
  m_axi_edge_list_ptr_ARLEN,
  m_axi_edge_list_ptr_ARLOCK,
  m_axi_edge_list_ptr_ARPROT,
  m_axi_edge_list_ptr_ARQOS,
  m_axi_edge_list_ptr_ARREADY,
  m_axi_edge_list_ptr_ARSIZE,
  m_axi_edge_list_ptr_ARVALID,
  m_axi_edge_list_ptr_AWADDR,
  m_axi_edge_list_ptr_AWBURST,
  m_axi_edge_list_ptr_AWCACHE,
  m_axi_edge_list_ptr_AWID,
  m_axi_edge_list_ptr_AWLEN,
  m_axi_edge_list_ptr_AWLOCK,
  m_axi_edge_list_ptr_AWPROT,
  m_axi_edge_list_ptr_AWQOS,
  m_axi_edge_list_ptr_AWREADY,
  m_axi_edge_list_ptr_AWSIZE,
  m_axi_edge_list_ptr_AWVALID,
  m_axi_edge_list_ptr_BID,
  m_axi_edge_list_ptr_BREADY,
  m_axi_edge_list_ptr_BRESP,
  m_axi_edge_list_ptr_BVALID,
  m_axi_edge_list_ptr_RDATA,
  m_axi_edge_list_ptr_RID,
  m_axi_edge_list_ptr_RLAST,
  m_axi_edge_list_ptr_RREADY,
  m_axi_edge_list_ptr_RRESP,
  m_axi_edge_list_ptr_RVALID,
  m_axi_edge_list_ptr_WDATA,
  m_axi_edge_list_ptr_WLAST,
  m_axi_edge_list_ptr_WREADY,
  m_axi_edge_list_ptr_WSTRB,
  m_axi_edge_list_ptr_WVALID,
  m_axi_mat_C_ch_0_ARADDR,
  m_axi_mat_C_ch_0_ARBURST,
  m_axi_mat_C_ch_0_ARCACHE,
  m_axi_mat_C_ch_0_ARID,
  m_axi_mat_C_ch_0_ARLEN,
  m_axi_mat_C_ch_0_ARLOCK,
  m_axi_mat_C_ch_0_ARPROT,
  m_axi_mat_C_ch_0_ARQOS,
  m_axi_mat_C_ch_0_ARREADY,
  m_axi_mat_C_ch_0_ARSIZE,
  m_axi_mat_C_ch_0_ARVALID,
  m_axi_mat_C_ch_0_AWADDR,
  m_axi_mat_C_ch_0_AWBURST,
  m_axi_mat_C_ch_0_AWCACHE,
  m_axi_mat_C_ch_0_AWID,
  m_axi_mat_C_ch_0_AWLEN,
  m_axi_mat_C_ch_0_AWLOCK,
  m_axi_mat_C_ch_0_AWPROT,
  m_axi_mat_C_ch_0_AWQOS,
  m_axi_mat_C_ch_0_AWREADY,
  m_axi_mat_C_ch_0_AWSIZE,
  m_axi_mat_C_ch_0_AWVALID,
  m_axi_mat_C_ch_0_BID,
  m_axi_mat_C_ch_0_BREADY,
  m_axi_mat_C_ch_0_BRESP,
  m_axi_mat_C_ch_0_BVALID,
  m_axi_mat_C_ch_0_RDATA,
  m_axi_mat_C_ch_0_RID,
  m_axi_mat_C_ch_0_RLAST,
  m_axi_mat_C_ch_0_RREADY,
  m_axi_mat_C_ch_0_RRESP,
  m_axi_mat_C_ch_0_RVALID,
  m_axi_mat_C_ch_0_WDATA,
  m_axi_mat_C_ch_0_WLAST,
  m_axi_mat_C_ch_0_WREADY,
  m_axi_mat_C_ch_0_WSTRB,
  m_axi_mat_C_ch_0_WVALID,
  m_axi_mat_C_ch_1_ARADDR,
  m_axi_mat_C_ch_1_ARBURST,
  m_axi_mat_C_ch_1_ARCACHE,
  m_axi_mat_C_ch_1_ARID,
  m_axi_mat_C_ch_1_ARLEN,
  m_axi_mat_C_ch_1_ARLOCK,
  m_axi_mat_C_ch_1_ARPROT,
  m_axi_mat_C_ch_1_ARQOS,
  m_axi_mat_C_ch_1_ARREADY,
  m_axi_mat_C_ch_1_ARSIZE,
  m_axi_mat_C_ch_1_ARVALID,
  m_axi_mat_C_ch_1_AWADDR,
  m_axi_mat_C_ch_1_AWBURST,
  m_axi_mat_C_ch_1_AWCACHE,
  m_axi_mat_C_ch_1_AWID,
  m_axi_mat_C_ch_1_AWLEN,
  m_axi_mat_C_ch_1_AWLOCK,
  m_axi_mat_C_ch_1_AWPROT,
  m_axi_mat_C_ch_1_AWQOS,
  m_axi_mat_C_ch_1_AWREADY,
  m_axi_mat_C_ch_1_AWSIZE,
  m_axi_mat_C_ch_1_AWVALID,
  m_axi_mat_C_ch_1_BID,
  m_axi_mat_C_ch_1_BREADY,
  m_axi_mat_C_ch_1_BRESP,
  m_axi_mat_C_ch_1_BVALID,
  m_axi_mat_C_ch_1_RDATA,
  m_axi_mat_C_ch_1_RID,
  m_axi_mat_C_ch_1_RLAST,
  m_axi_mat_C_ch_1_RREADY,
  m_axi_mat_C_ch_1_RRESP,
  m_axi_mat_C_ch_1_RVALID,
  m_axi_mat_C_ch_1_WDATA,
  m_axi_mat_C_ch_1_WLAST,
  m_axi_mat_C_ch_1_WREADY,
  m_axi_mat_C_ch_1_WSTRB,
  m_axi_mat_C_ch_1_WVALID,
  m_axi_mat_C_ch_2_ARADDR,
  m_axi_mat_C_ch_2_ARBURST,
  m_axi_mat_C_ch_2_ARCACHE,
  m_axi_mat_C_ch_2_ARID,
  m_axi_mat_C_ch_2_ARLEN,
  m_axi_mat_C_ch_2_ARLOCK,
  m_axi_mat_C_ch_2_ARPROT,
  m_axi_mat_C_ch_2_ARQOS,
  m_axi_mat_C_ch_2_ARREADY,
  m_axi_mat_C_ch_2_ARSIZE,
  m_axi_mat_C_ch_2_ARVALID,
  m_axi_mat_C_ch_2_AWADDR,
  m_axi_mat_C_ch_2_AWBURST,
  m_axi_mat_C_ch_2_AWCACHE,
  m_axi_mat_C_ch_2_AWID,
  m_axi_mat_C_ch_2_AWLEN,
  m_axi_mat_C_ch_2_AWLOCK,
  m_axi_mat_C_ch_2_AWPROT,
  m_axi_mat_C_ch_2_AWQOS,
  m_axi_mat_C_ch_2_AWREADY,
  m_axi_mat_C_ch_2_AWSIZE,
  m_axi_mat_C_ch_2_AWVALID,
  m_axi_mat_C_ch_2_BID,
  m_axi_mat_C_ch_2_BREADY,
  m_axi_mat_C_ch_2_BRESP,
  m_axi_mat_C_ch_2_BVALID,
  m_axi_mat_C_ch_2_RDATA,
  m_axi_mat_C_ch_2_RID,
  m_axi_mat_C_ch_2_RLAST,
  m_axi_mat_C_ch_2_RREADY,
  m_axi_mat_C_ch_2_RRESP,
  m_axi_mat_C_ch_2_RVALID,
  m_axi_mat_C_ch_2_WDATA,
  m_axi_mat_C_ch_2_WLAST,
  m_axi_mat_C_ch_2_WREADY,
  m_axi_mat_C_ch_2_WSTRB,
  m_axi_mat_C_ch_2_WVALID,
  m_axi_mat_C_ch_3_ARADDR,
  m_axi_mat_C_ch_3_ARBURST,
  m_axi_mat_C_ch_3_ARCACHE,
  m_axi_mat_C_ch_3_ARID,
  m_axi_mat_C_ch_3_ARLEN,
  m_axi_mat_C_ch_3_ARLOCK,
  m_axi_mat_C_ch_3_ARPROT,
  m_axi_mat_C_ch_3_ARQOS,
  m_axi_mat_C_ch_3_ARREADY,
  m_axi_mat_C_ch_3_ARSIZE,
  m_axi_mat_C_ch_3_ARVALID,
  m_axi_mat_C_ch_3_AWADDR,
  m_axi_mat_C_ch_3_AWBURST,
  m_axi_mat_C_ch_3_AWCACHE,
  m_axi_mat_C_ch_3_AWID,
  m_axi_mat_C_ch_3_AWLEN,
  m_axi_mat_C_ch_3_AWLOCK,
  m_axi_mat_C_ch_3_AWPROT,
  m_axi_mat_C_ch_3_AWQOS,
  m_axi_mat_C_ch_3_AWREADY,
  m_axi_mat_C_ch_3_AWSIZE,
  m_axi_mat_C_ch_3_AWVALID,
  m_axi_mat_C_ch_3_BID,
  m_axi_mat_C_ch_3_BREADY,
  m_axi_mat_C_ch_3_BRESP,
  m_axi_mat_C_ch_3_BVALID,
  m_axi_mat_C_ch_3_RDATA,
  m_axi_mat_C_ch_3_RID,
  m_axi_mat_C_ch_3_RLAST,
  m_axi_mat_C_ch_3_RREADY,
  m_axi_mat_C_ch_3_RRESP,
  m_axi_mat_C_ch_3_RVALID,
  m_axi_mat_C_ch_3_WDATA,
  m_axi_mat_C_ch_3_WLAST,
  m_axi_mat_C_ch_3_WREADY,
  m_axi_mat_C_ch_3_WSTRB,
  m_axi_mat_C_ch_3_WVALID,
  m_axi_mat_C_ch_4_ARADDR,
  m_axi_mat_C_ch_4_ARBURST,
  m_axi_mat_C_ch_4_ARCACHE,
  m_axi_mat_C_ch_4_ARID,
  m_axi_mat_C_ch_4_ARLEN,
  m_axi_mat_C_ch_4_ARLOCK,
  m_axi_mat_C_ch_4_ARPROT,
  m_axi_mat_C_ch_4_ARQOS,
  m_axi_mat_C_ch_4_ARREADY,
  m_axi_mat_C_ch_4_ARSIZE,
  m_axi_mat_C_ch_4_ARVALID,
  m_axi_mat_C_ch_4_AWADDR,
  m_axi_mat_C_ch_4_AWBURST,
  m_axi_mat_C_ch_4_AWCACHE,
  m_axi_mat_C_ch_4_AWID,
  m_axi_mat_C_ch_4_AWLEN,
  m_axi_mat_C_ch_4_AWLOCK,
  m_axi_mat_C_ch_4_AWPROT,
  m_axi_mat_C_ch_4_AWQOS,
  m_axi_mat_C_ch_4_AWREADY,
  m_axi_mat_C_ch_4_AWSIZE,
  m_axi_mat_C_ch_4_AWVALID,
  m_axi_mat_C_ch_4_BID,
  m_axi_mat_C_ch_4_BREADY,
  m_axi_mat_C_ch_4_BRESP,
  m_axi_mat_C_ch_4_BVALID,
  m_axi_mat_C_ch_4_RDATA,
  m_axi_mat_C_ch_4_RID,
  m_axi_mat_C_ch_4_RLAST,
  m_axi_mat_C_ch_4_RREADY,
  m_axi_mat_C_ch_4_RRESP,
  m_axi_mat_C_ch_4_RVALID,
  m_axi_mat_C_ch_4_WDATA,
  m_axi_mat_C_ch_4_WLAST,
  m_axi_mat_C_ch_4_WREADY,
  m_axi_mat_C_ch_4_WSTRB,
  m_axi_mat_C_ch_4_WVALID,
  m_axi_mat_C_ch_5_ARADDR,
  m_axi_mat_C_ch_5_ARBURST,
  m_axi_mat_C_ch_5_ARCACHE,
  m_axi_mat_C_ch_5_ARID,
  m_axi_mat_C_ch_5_ARLEN,
  m_axi_mat_C_ch_5_ARLOCK,
  m_axi_mat_C_ch_5_ARPROT,
  m_axi_mat_C_ch_5_ARQOS,
  m_axi_mat_C_ch_5_ARREADY,
  m_axi_mat_C_ch_5_ARSIZE,
  m_axi_mat_C_ch_5_ARVALID,
  m_axi_mat_C_ch_5_AWADDR,
  m_axi_mat_C_ch_5_AWBURST,
  m_axi_mat_C_ch_5_AWCACHE,
  m_axi_mat_C_ch_5_AWID,
  m_axi_mat_C_ch_5_AWLEN,
  m_axi_mat_C_ch_5_AWLOCK,
  m_axi_mat_C_ch_5_AWPROT,
  m_axi_mat_C_ch_5_AWQOS,
  m_axi_mat_C_ch_5_AWREADY,
  m_axi_mat_C_ch_5_AWSIZE,
  m_axi_mat_C_ch_5_AWVALID,
  m_axi_mat_C_ch_5_BID,
  m_axi_mat_C_ch_5_BREADY,
  m_axi_mat_C_ch_5_BRESP,
  m_axi_mat_C_ch_5_BVALID,
  m_axi_mat_C_ch_5_RDATA,
  m_axi_mat_C_ch_5_RID,
  m_axi_mat_C_ch_5_RLAST,
  m_axi_mat_C_ch_5_RREADY,
  m_axi_mat_C_ch_5_RRESP,
  m_axi_mat_C_ch_5_RVALID,
  m_axi_mat_C_ch_5_WDATA,
  m_axi_mat_C_ch_5_WLAST,
  m_axi_mat_C_ch_5_WREADY,
  m_axi_mat_C_ch_5_WSTRB,
  m_axi_mat_C_ch_5_WVALID,
  m_axi_mat_C_ch_6_ARADDR,
  m_axi_mat_C_ch_6_ARBURST,
  m_axi_mat_C_ch_6_ARCACHE,
  m_axi_mat_C_ch_6_ARID,
  m_axi_mat_C_ch_6_ARLEN,
  m_axi_mat_C_ch_6_ARLOCK,
  m_axi_mat_C_ch_6_ARPROT,
  m_axi_mat_C_ch_6_ARQOS,
  m_axi_mat_C_ch_6_ARREADY,
  m_axi_mat_C_ch_6_ARSIZE,
  m_axi_mat_C_ch_6_ARVALID,
  m_axi_mat_C_ch_6_AWADDR,
  m_axi_mat_C_ch_6_AWBURST,
  m_axi_mat_C_ch_6_AWCACHE,
  m_axi_mat_C_ch_6_AWID,
  m_axi_mat_C_ch_6_AWLEN,
  m_axi_mat_C_ch_6_AWLOCK,
  m_axi_mat_C_ch_6_AWPROT,
  m_axi_mat_C_ch_6_AWQOS,
  m_axi_mat_C_ch_6_AWREADY,
  m_axi_mat_C_ch_6_AWSIZE,
  m_axi_mat_C_ch_6_AWVALID,
  m_axi_mat_C_ch_6_BID,
  m_axi_mat_C_ch_6_BREADY,
  m_axi_mat_C_ch_6_BRESP,
  m_axi_mat_C_ch_6_BVALID,
  m_axi_mat_C_ch_6_RDATA,
  m_axi_mat_C_ch_6_RID,
  m_axi_mat_C_ch_6_RLAST,
  m_axi_mat_C_ch_6_RREADY,
  m_axi_mat_C_ch_6_RRESP,
  m_axi_mat_C_ch_6_RVALID,
  m_axi_mat_C_ch_6_WDATA,
  m_axi_mat_C_ch_6_WLAST,
  m_axi_mat_C_ch_6_WREADY,
  m_axi_mat_C_ch_6_WSTRB,
  m_axi_mat_C_ch_6_WVALID,
  m_axi_mat_C_ch_7_ARADDR,
  m_axi_mat_C_ch_7_ARBURST,
  m_axi_mat_C_ch_7_ARCACHE,
  m_axi_mat_C_ch_7_ARID,
  m_axi_mat_C_ch_7_ARLEN,
  m_axi_mat_C_ch_7_ARLOCK,
  m_axi_mat_C_ch_7_ARPROT,
  m_axi_mat_C_ch_7_ARQOS,
  m_axi_mat_C_ch_7_ARREADY,
  m_axi_mat_C_ch_7_ARSIZE,
  m_axi_mat_C_ch_7_ARVALID,
  m_axi_mat_C_ch_7_AWADDR,
  m_axi_mat_C_ch_7_AWBURST,
  m_axi_mat_C_ch_7_AWCACHE,
  m_axi_mat_C_ch_7_AWID,
  m_axi_mat_C_ch_7_AWLEN,
  m_axi_mat_C_ch_7_AWLOCK,
  m_axi_mat_C_ch_7_AWPROT,
  m_axi_mat_C_ch_7_AWQOS,
  m_axi_mat_C_ch_7_AWREADY,
  m_axi_mat_C_ch_7_AWSIZE,
  m_axi_mat_C_ch_7_AWVALID,
  m_axi_mat_C_ch_7_BID,
  m_axi_mat_C_ch_7_BREADY,
  m_axi_mat_C_ch_7_BRESP,
  m_axi_mat_C_ch_7_BVALID,
  m_axi_mat_C_ch_7_RDATA,
  m_axi_mat_C_ch_7_RID,
  m_axi_mat_C_ch_7_RLAST,
  m_axi_mat_C_ch_7_RREADY,
  m_axi_mat_C_ch_7_RRESP,
  m_axi_mat_C_ch_7_RVALID,
  m_axi_mat_C_ch_7_WDATA,
  m_axi_mat_C_ch_7_WLAST,
  m_axi_mat_C_ch_7_WREADY,
  m_axi_mat_C_ch_7_WSTRB,
  m_axi_mat_C_ch_7_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 9;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  (* RS_HS = "s_axi_control_AW.valid" *)input s_axi_control_AWVALID;
  (* RS_HS = "s_axi_control_AW.ready" *)output s_axi_control_AWREADY;
  (* RS_HS = "s_axi_control_AW.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  (* RS_HS = "s_axi_control_W.valid" *)input s_axi_control_WVALID;
  (* RS_HS = "s_axi_control_W.ready" *)output s_axi_control_WREADY;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  (* RS_HS = "s_axi_control_AR.valid" *)input s_axi_control_ARVALID;
  (* RS_HS = "s_axi_control_AR.ready" *)output s_axi_control_ARREADY;
  (* RS_HS = "s_axi_control_AR.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  (* RS_HS = "s_axi_control_R.valid" *)output s_axi_control_RVALID;
  (* RS_HS = "s_axi_control_R.ready" *)input s_axi_control_RREADY;
  (* RS_HS = "s_axi_control_R.data" *)output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  (* RS_HS = "s_axi_control_R.data" *)output [1:0] s_axi_control_RRESP;
  (* RS_HS = "s_axi_control_B.valid" *)output s_axi_control_BVALID;
  (* RS_HS = "s_axi_control_B.ready" *)input s_axi_control_BREADY;
  (* RS_HS = "s_axi_control_B.data" *)output [1:0] s_axi_control_BRESP;
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_FF = "interrupt" *)output interrupt;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [63:0] m_axi_edge_list_ch_0_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [1:0] m_axi_edge_list_ch_0_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [3:0] m_axi_edge_list_ch_0_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [0:0] m_axi_edge_list_ch_0_ARID;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [7:0] m_axi_edge_list_ch_0_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output m_axi_edge_list_ch_0_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [2:0] m_axi_edge_list_ch_0_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [3:0] m_axi_edge_list_ch_0_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.ready" *)input m_axi_edge_list_ch_0_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.data" *)output [2:0] m_axi_edge_list_ch_0_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_0_AR.valid" *)output m_axi_edge_list_ch_0_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [63:0] m_axi_edge_list_ch_0_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [1:0] m_axi_edge_list_ch_0_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [3:0] m_axi_edge_list_ch_0_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [0:0] m_axi_edge_list_ch_0_AWID;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [7:0] m_axi_edge_list_ch_0_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output m_axi_edge_list_ch_0_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [2:0] m_axi_edge_list_ch_0_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [3:0] m_axi_edge_list_ch_0_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.ready" *)input m_axi_edge_list_ch_0_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.data" *)output [2:0] m_axi_edge_list_ch_0_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_0_AW.valid" *)output m_axi_edge_list_ch_0_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_0_B.data" *)input [0:0] m_axi_edge_list_ch_0_BID;
  (* RS_HS = "m_axi_edge_list_ch_0_B.ready" *)output m_axi_edge_list_ch_0_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_0_B.data" *)input [1:0] m_axi_edge_list_ch_0_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_0_B.valid" *)input m_axi_edge_list_ch_0_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_0_R.data" *)input [511:0] m_axi_edge_list_ch_0_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_0_R.data" *)input [0:0] m_axi_edge_list_ch_0_RID;
  (* RS_HS = "m_axi_edge_list_ch_0_R.data" *)input m_axi_edge_list_ch_0_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_0_R.ready" *)output m_axi_edge_list_ch_0_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_0_R.data" *)input [1:0] m_axi_edge_list_ch_0_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_0_R.valid" *)input m_axi_edge_list_ch_0_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_0_W.data" *)output [511:0] m_axi_edge_list_ch_0_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_0_W.data" *)output m_axi_edge_list_ch_0_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_0_W.ready" *)input m_axi_edge_list_ch_0_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_0_W.data" *)output [63:0] m_axi_edge_list_ch_0_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_0_W.valid" *)output m_axi_edge_list_ch_0_WVALID;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [63:0] m_axi_edge_list_ch_1_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [1:0] m_axi_edge_list_ch_1_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [3:0] m_axi_edge_list_ch_1_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [0:0] m_axi_edge_list_ch_1_ARID;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [7:0] m_axi_edge_list_ch_1_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output m_axi_edge_list_ch_1_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [2:0] m_axi_edge_list_ch_1_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [3:0] m_axi_edge_list_ch_1_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.ready" *)input m_axi_edge_list_ch_1_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.data" *)output [2:0] m_axi_edge_list_ch_1_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_1_AR.valid" *)output m_axi_edge_list_ch_1_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [63:0] m_axi_edge_list_ch_1_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [1:0] m_axi_edge_list_ch_1_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [3:0] m_axi_edge_list_ch_1_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [0:0] m_axi_edge_list_ch_1_AWID;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [7:0] m_axi_edge_list_ch_1_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output m_axi_edge_list_ch_1_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [2:0] m_axi_edge_list_ch_1_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [3:0] m_axi_edge_list_ch_1_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.ready" *)input m_axi_edge_list_ch_1_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.data" *)output [2:0] m_axi_edge_list_ch_1_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_1_AW.valid" *)output m_axi_edge_list_ch_1_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_1_B.data" *)input [0:0] m_axi_edge_list_ch_1_BID;
  (* RS_HS = "m_axi_edge_list_ch_1_B.ready" *)output m_axi_edge_list_ch_1_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_1_B.data" *)input [1:0] m_axi_edge_list_ch_1_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_1_B.valid" *)input m_axi_edge_list_ch_1_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_1_R.data" *)input [511:0] m_axi_edge_list_ch_1_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_1_R.data" *)input [0:0] m_axi_edge_list_ch_1_RID;
  (* RS_HS = "m_axi_edge_list_ch_1_R.data" *)input m_axi_edge_list_ch_1_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_1_R.ready" *)output m_axi_edge_list_ch_1_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_1_R.data" *)input [1:0] m_axi_edge_list_ch_1_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_1_R.valid" *)input m_axi_edge_list_ch_1_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_1_W.data" *)output [511:0] m_axi_edge_list_ch_1_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_1_W.data" *)output m_axi_edge_list_ch_1_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_1_W.ready" *)input m_axi_edge_list_ch_1_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_1_W.data" *)output [63:0] m_axi_edge_list_ch_1_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_1_W.valid" *)output m_axi_edge_list_ch_1_WVALID;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [63:0] m_axi_edge_list_ch_2_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [1:0] m_axi_edge_list_ch_2_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [3:0] m_axi_edge_list_ch_2_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [0:0] m_axi_edge_list_ch_2_ARID;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [7:0] m_axi_edge_list_ch_2_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output m_axi_edge_list_ch_2_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [2:0] m_axi_edge_list_ch_2_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [3:0] m_axi_edge_list_ch_2_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.ready" *)input m_axi_edge_list_ch_2_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.data" *)output [2:0] m_axi_edge_list_ch_2_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_2_AR.valid" *)output m_axi_edge_list_ch_2_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [63:0] m_axi_edge_list_ch_2_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [1:0] m_axi_edge_list_ch_2_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [3:0] m_axi_edge_list_ch_2_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [0:0] m_axi_edge_list_ch_2_AWID;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [7:0] m_axi_edge_list_ch_2_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output m_axi_edge_list_ch_2_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [2:0] m_axi_edge_list_ch_2_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [3:0] m_axi_edge_list_ch_2_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.ready" *)input m_axi_edge_list_ch_2_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.data" *)output [2:0] m_axi_edge_list_ch_2_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_2_AW.valid" *)output m_axi_edge_list_ch_2_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_2_B.data" *)input [0:0] m_axi_edge_list_ch_2_BID;
  (* RS_HS = "m_axi_edge_list_ch_2_B.ready" *)output m_axi_edge_list_ch_2_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_2_B.data" *)input [1:0] m_axi_edge_list_ch_2_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_2_B.valid" *)input m_axi_edge_list_ch_2_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_2_R.data" *)input [511:0] m_axi_edge_list_ch_2_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_2_R.data" *)input [0:0] m_axi_edge_list_ch_2_RID;
  (* RS_HS = "m_axi_edge_list_ch_2_R.data" *)input m_axi_edge_list_ch_2_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_2_R.ready" *)output m_axi_edge_list_ch_2_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_2_R.data" *)input [1:0] m_axi_edge_list_ch_2_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_2_R.valid" *)input m_axi_edge_list_ch_2_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_2_W.data" *)output [511:0] m_axi_edge_list_ch_2_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_2_W.data" *)output m_axi_edge_list_ch_2_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_2_W.ready" *)input m_axi_edge_list_ch_2_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_2_W.data" *)output [63:0] m_axi_edge_list_ch_2_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_2_W.valid" *)output m_axi_edge_list_ch_2_WVALID;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [63:0] m_axi_edge_list_ch_3_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [1:0] m_axi_edge_list_ch_3_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [3:0] m_axi_edge_list_ch_3_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [0:0] m_axi_edge_list_ch_3_ARID;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [7:0] m_axi_edge_list_ch_3_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output m_axi_edge_list_ch_3_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [2:0] m_axi_edge_list_ch_3_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [3:0] m_axi_edge_list_ch_3_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.ready" *)input m_axi_edge_list_ch_3_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.data" *)output [2:0] m_axi_edge_list_ch_3_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_3_AR.valid" *)output m_axi_edge_list_ch_3_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [63:0] m_axi_edge_list_ch_3_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [1:0] m_axi_edge_list_ch_3_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [3:0] m_axi_edge_list_ch_3_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [0:0] m_axi_edge_list_ch_3_AWID;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [7:0] m_axi_edge_list_ch_3_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output m_axi_edge_list_ch_3_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [2:0] m_axi_edge_list_ch_3_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [3:0] m_axi_edge_list_ch_3_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.ready" *)input m_axi_edge_list_ch_3_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.data" *)output [2:0] m_axi_edge_list_ch_3_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_3_AW.valid" *)output m_axi_edge_list_ch_3_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_3_B.data" *)input [0:0] m_axi_edge_list_ch_3_BID;
  (* RS_HS = "m_axi_edge_list_ch_3_B.ready" *)output m_axi_edge_list_ch_3_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_3_B.data" *)input [1:0] m_axi_edge_list_ch_3_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_3_B.valid" *)input m_axi_edge_list_ch_3_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_3_R.data" *)input [511:0] m_axi_edge_list_ch_3_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_3_R.data" *)input [0:0] m_axi_edge_list_ch_3_RID;
  (* RS_HS = "m_axi_edge_list_ch_3_R.data" *)input m_axi_edge_list_ch_3_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_3_R.ready" *)output m_axi_edge_list_ch_3_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_3_R.data" *)input [1:0] m_axi_edge_list_ch_3_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_3_R.valid" *)input m_axi_edge_list_ch_3_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_3_W.data" *)output [511:0] m_axi_edge_list_ch_3_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_3_W.data" *)output m_axi_edge_list_ch_3_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_3_W.ready" *)input m_axi_edge_list_ch_3_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_3_W.data" *)output [63:0] m_axi_edge_list_ch_3_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_3_W.valid" *)output m_axi_edge_list_ch_3_WVALID;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [63:0] m_axi_edge_list_ch_4_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [1:0] m_axi_edge_list_ch_4_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [3:0] m_axi_edge_list_ch_4_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [0:0] m_axi_edge_list_ch_4_ARID;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [7:0] m_axi_edge_list_ch_4_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output m_axi_edge_list_ch_4_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [2:0] m_axi_edge_list_ch_4_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [3:0] m_axi_edge_list_ch_4_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.ready" *)input m_axi_edge_list_ch_4_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.data" *)output [2:0] m_axi_edge_list_ch_4_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_4_AR.valid" *)output m_axi_edge_list_ch_4_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [63:0] m_axi_edge_list_ch_4_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [1:0] m_axi_edge_list_ch_4_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [3:0] m_axi_edge_list_ch_4_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [0:0] m_axi_edge_list_ch_4_AWID;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [7:0] m_axi_edge_list_ch_4_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output m_axi_edge_list_ch_4_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [2:0] m_axi_edge_list_ch_4_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [3:0] m_axi_edge_list_ch_4_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.ready" *)input m_axi_edge_list_ch_4_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.data" *)output [2:0] m_axi_edge_list_ch_4_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_4_AW.valid" *)output m_axi_edge_list_ch_4_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_4_B.data" *)input [0:0] m_axi_edge_list_ch_4_BID;
  (* RS_HS = "m_axi_edge_list_ch_4_B.ready" *)output m_axi_edge_list_ch_4_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_4_B.data" *)input [1:0] m_axi_edge_list_ch_4_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_4_B.valid" *)input m_axi_edge_list_ch_4_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_4_R.data" *)input [511:0] m_axi_edge_list_ch_4_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_4_R.data" *)input [0:0] m_axi_edge_list_ch_4_RID;
  (* RS_HS = "m_axi_edge_list_ch_4_R.data" *)input m_axi_edge_list_ch_4_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_4_R.ready" *)output m_axi_edge_list_ch_4_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_4_R.data" *)input [1:0] m_axi_edge_list_ch_4_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_4_R.valid" *)input m_axi_edge_list_ch_4_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_4_W.data" *)output [511:0] m_axi_edge_list_ch_4_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_4_W.data" *)output m_axi_edge_list_ch_4_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_4_W.ready" *)input m_axi_edge_list_ch_4_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_4_W.data" *)output [63:0] m_axi_edge_list_ch_4_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_4_W.valid" *)output m_axi_edge_list_ch_4_WVALID;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [63:0] m_axi_edge_list_ch_5_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [1:0] m_axi_edge_list_ch_5_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [3:0] m_axi_edge_list_ch_5_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [0:0] m_axi_edge_list_ch_5_ARID;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [7:0] m_axi_edge_list_ch_5_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output m_axi_edge_list_ch_5_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [2:0] m_axi_edge_list_ch_5_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [3:0] m_axi_edge_list_ch_5_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.ready" *)input m_axi_edge_list_ch_5_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.data" *)output [2:0] m_axi_edge_list_ch_5_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_5_AR.valid" *)output m_axi_edge_list_ch_5_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [63:0] m_axi_edge_list_ch_5_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [1:0] m_axi_edge_list_ch_5_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [3:0] m_axi_edge_list_ch_5_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [0:0] m_axi_edge_list_ch_5_AWID;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [7:0] m_axi_edge_list_ch_5_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output m_axi_edge_list_ch_5_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [2:0] m_axi_edge_list_ch_5_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [3:0] m_axi_edge_list_ch_5_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.ready" *)input m_axi_edge_list_ch_5_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.data" *)output [2:0] m_axi_edge_list_ch_5_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_5_AW.valid" *)output m_axi_edge_list_ch_5_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_5_B.data" *)input [0:0] m_axi_edge_list_ch_5_BID;
  (* RS_HS = "m_axi_edge_list_ch_5_B.ready" *)output m_axi_edge_list_ch_5_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_5_B.data" *)input [1:0] m_axi_edge_list_ch_5_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_5_B.valid" *)input m_axi_edge_list_ch_5_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_5_R.data" *)input [511:0] m_axi_edge_list_ch_5_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_5_R.data" *)input [0:0] m_axi_edge_list_ch_5_RID;
  (* RS_HS = "m_axi_edge_list_ch_5_R.data" *)input m_axi_edge_list_ch_5_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_5_R.ready" *)output m_axi_edge_list_ch_5_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_5_R.data" *)input [1:0] m_axi_edge_list_ch_5_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_5_R.valid" *)input m_axi_edge_list_ch_5_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_5_W.data" *)output [511:0] m_axi_edge_list_ch_5_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_5_W.data" *)output m_axi_edge_list_ch_5_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_5_W.ready" *)input m_axi_edge_list_ch_5_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_5_W.data" *)output [63:0] m_axi_edge_list_ch_5_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_5_W.valid" *)output m_axi_edge_list_ch_5_WVALID;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [63:0] m_axi_edge_list_ch_6_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [1:0] m_axi_edge_list_ch_6_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [3:0] m_axi_edge_list_ch_6_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [0:0] m_axi_edge_list_ch_6_ARID;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [7:0] m_axi_edge_list_ch_6_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output m_axi_edge_list_ch_6_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [2:0] m_axi_edge_list_ch_6_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [3:0] m_axi_edge_list_ch_6_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.ready" *)input m_axi_edge_list_ch_6_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.data" *)output [2:0] m_axi_edge_list_ch_6_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_6_AR.valid" *)output m_axi_edge_list_ch_6_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [63:0] m_axi_edge_list_ch_6_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [1:0] m_axi_edge_list_ch_6_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [3:0] m_axi_edge_list_ch_6_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [0:0] m_axi_edge_list_ch_6_AWID;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [7:0] m_axi_edge_list_ch_6_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output m_axi_edge_list_ch_6_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [2:0] m_axi_edge_list_ch_6_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [3:0] m_axi_edge_list_ch_6_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.ready" *)input m_axi_edge_list_ch_6_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.data" *)output [2:0] m_axi_edge_list_ch_6_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_6_AW.valid" *)output m_axi_edge_list_ch_6_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_6_B.data" *)input [0:0] m_axi_edge_list_ch_6_BID;
  (* RS_HS = "m_axi_edge_list_ch_6_B.ready" *)output m_axi_edge_list_ch_6_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_6_B.data" *)input [1:0] m_axi_edge_list_ch_6_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_6_B.valid" *)input m_axi_edge_list_ch_6_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_6_R.data" *)input [511:0] m_axi_edge_list_ch_6_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_6_R.data" *)input [0:0] m_axi_edge_list_ch_6_RID;
  (* RS_HS = "m_axi_edge_list_ch_6_R.data" *)input m_axi_edge_list_ch_6_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_6_R.ready" *)output m_axi_edge_list_ch_6_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_6_R.data" *)input [1:0] m_axi_edge_list_ch_6_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_6_R.valid" *)input m_axi_edge_list_ch_6_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_6_W.data" *)output [511:0] m_axi_edge_list_ch_6_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_6_W.data" *)output m_axi_edge_list_ch_6_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_6_W.ready" *)input m_axi_edge_list_ch_6_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_6_W.data" *)output [63:0] m_axi_edge_list_ch_6_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_6_W.valid" *)output m_axi_edge_list_ch_6_WVALID;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [63:0] m_axi_edge_list_ch_7_ARADDR;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [1:0] m_axi_edge_list_ch_7_ARBURST;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [3:0] m_axi_edge_list_ch_7_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [0:0] m_axi_edge_list_ch_7_ARID;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [7:0] m_axi_edge_list_ch_7_ARLEN;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output m_axi_edge_list_ch_7_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [2:0] m_axi_edge_list_ch_7_ARPROT;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [3:0] m_axi_edge_list_ch_7_ARQOS;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.ready" *)input m_axi_edge_list_ch_7_ARREADY;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.data" *)output [2:0] m_axi_edge_list_ch_7_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ch_7_AR.valid" *)output m_axi_edge_list_ch_7_ARVALID;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [63:0] m_axi_edge_list_ch_7_AWADDR;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [1:0] m_axi_edge_list_ch_7_AWBURST;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [3:0] m_axi_edge_list_ch_7_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [0:0] m_axi_edge_list_ch_7_AWID;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [7:0] m_axi_edge_list_ch_7_AWLEN;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output m_axi_edge_list_ch_7_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [2:0] m_axi_edge_list_ch_7_AWPROT;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [3:0] m_axi_edge_list_ch_7_AWQOS;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.ready" *)input m_axi_edge_list_ch_7_AWREADY;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.data" *)output [2:0] m_axi_edge_list_ch_7_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ch_7_AW.valid" *)output m_axi_edge_list_ch_7_AWVALID;
  (* RS_HS = "m_axi_edge_list_ch_7_B.data" *)input [0:0] m_axi_edge_list_ch_7_BID;
  (* RS_HS = "m_axi_edge_list_ch_7_B.ready" *)output m_axi_edge_list_ch_7_BREADY;
  (* RS_HS = "m_axi_edge_list_ch_7_B.data" *)input [1:0] m_axi_edge_list_ch_7_BRESP;
  (* RS_HS = "m_axi_edge_list_ch_7_B.valid" *)input m_axi_edge_list_ch_7_BVALID;
  (* RS_HS = "m_axi_edge_list_ch_7_R.data" *)input [511:0] m_axi_edge_list_ch_7_RDATA;
  (* RS_HS = "m_axi_edge_list_ch_7_R.data" *)input [0:0] m_axi_edge_list_ch_7_RID;
  (* RS_HS = "m_axi_edge_list_ch_7_R.data" *)input m_axi_edge_list_ch_7_RLAST;
  (* RS_HS = "m_axi_edge_list_ch_7_R.ready" *)output m_axi_edge_list_ch_7_RREADY;
  (* RS_HS = "m_axi_edge_list_ch_7_R.data" *)input [1:0] m_axi_edge_list_ch_7_RRESP;
  (* RS_HS = "m_axi_edge_list_ch_7_R.valid" *)input m_axi_edge_list_ch_7_RVALID;
  (* RS_HS = "m_axi_edge_list_ch_7_W.data" *)output [511:0] m_axi_edge_list_ch_7_WDATA;
  (* RS_HS = "m_axi_edge_list_ch_7_W.data" *)output m_axi_edge_list_ch_7_WLAST;
  (* RS_HS = "m_axi_edge_list_ch_7_W.ready" *)input m_axi_edge_list_ch_7_WREADY;
  (* RS_HS = "m_axi_edge_list_ch_7_W.data" *)output [63:0] m_axi_edge_list_ch_7_WSTRB;
  (* RS_HS = "m_axi_edge_list_ch_7_W.valid" *)output m_axi_edge_list_ch_7_WVALID;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [63:0] m_axi_mat_B_ch_0_ARADDR;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [1:0] m_axi_mat_B_ch_0_ARBURST;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [3:0] m_axi_mat_B_ch_0_ARCACHE;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [0:0] m_axi_mat_B_ch_0_ARID;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [7:0] m_axi_mat_B_ch_0_ARLEN;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output m_axi_mat_B_ch_0_ARLOCK;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [2:0] m_axi_mat_B_ch_0_ARPROT;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [3:0] m_axi_mat_B_ch_0_ARQOS;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.ready" *)input m_axi_mat_B_ch_0_ARREADY;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.data" *)output [2:0] m_axi_mat_B_ch_0_ARSIZE;
  (* RS_HS = "m_axi_mat_B_ch_0_AR.valid" *)output m_axi_mat_B_ch_0_ARVALID;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [63:0] m_axi_mat_B_ch_0_AWADDR;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [1:0] m_axi_mat_B_ch_0_AWBURST;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [3:0] m_axi_mat_B_ch_0_AWCACHE;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [0:0] m_axi_mat_B_ch_0_AWID;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [7:0] m_axi_mat_B_ch_0_AWLEN;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output m_axi_mat_B_ch_0_AWLOCK;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [2:0] m_axi_mat_B_ch_0_AWPROT;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [3:0] m_axi_mat_B_ch_0_AWQOS;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.ready" *)input m_axi_mat_B_ch_0_AWREADY;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.data" *)output [2:0] m_axi_mat_B_ch_0_AWSIZE;
  (* RS_HS = "m_axi_mat_B_ch_0_AW.valid" *)output m_axi_mat_B_ch_0_AWVALID;
  (* RS_HS = "m_axi_mat_B_ch_0_B.data" *)input [0:0] m_axi_mat_B_ch_0_BID;
  (* RS_HS = "m_axi_mat_B_ch_0_B.ready" *)output m_axi_mat_B_ch_0_BREADY;
  (* RS_HS = "m_axi_mat_B_ch_0_B.data" *)input [1:0] m_axi_mat_B_ch_0_BRESP;
  (* RS_HS = "m_axi_mat_B_ch_0_B.valid" *)input m_axi_mat_B_ch_0_BVALID;
  (* RS_HS = "m_axi_mat_B_ch_0_R.data" *)input [511:0] m_axi_mat_B_ch_0_RDATA;
  (* RS_HS = "m_axi_mat_B_ch_0_R.data" *)input [0:0] m_axi_mat_B_ch_0_RID;
  (* RS_HS = "m_axi_mat_B_ch_0_R.data" *)input m_axi_mat_B_ch_0_RLAST;
  (* RS_HS = "m_axi_mat_B_ch_0_R.ready" *)output m_axi_mat_B_ch_0_RREADY;
  (* RS_HS = "m_axi_mat_B_ch_0_R.data" *)input [1:0] m_axi_mat_B_ch_0_RRESP;
  (* RS_HS = "m_axi_mat_B_ch_0_R.valid" *)input m_axi_mat_B_ch_0_RVALID;
  (* RS_HS = "m_axi_mat_B_ch_0_W.data" *)output [511:0] m_axi_mat_B_ch_0_WDATA;
  (* RS_HS = "m_axi_mat_B_ch_0_W.data" *)output m_axi_mat_B_ch_0_WLAST;
  (* RS_HS = "m_axi_mat_B_ch_0_W.ready" *)input m_axi_mat_B_ch_0_WREADY;
  (* RS_HS = "m_axi_mat_B_ch_0_W.data" *)output [63:0] m_axi_mat_B_ch_0_WSTRB;
  (* RS_HS = "m_axi_mat_B_ch_0_W.valid" *)output m_axi_mat_B_ch_0_WVALID;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [63:0] m_axi_mat_B_ch_1_ARADDR;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [1:0] m_axi_mat_B_ch_1_ARBURST;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [3:0] m_axi_mat_B_ch_1_ARCACHE;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [0:0] m_axi_mat_B_ch_1_ARID;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [7:0] m_axi_mat_B_ch_1_ARLEN;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output m_axi_mat_B_ch_1_ARLOCK;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [2:0] m_axi_mat_B_ch_1_ARPROT;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [3:0] m_axi_mat_B_ch_1_ARQOS;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.ready" *)input m_axi_mat_B_ch_1_ARREADY;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.data" *)output [2:0] m_axi_mat_B_ch_1_ARSIZE;
  (* RS_HS = "m_axi_mat_B_ch_1_AR.valid" *)output m_axi_mat_B_ch_1_ARVALID;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [63:0] m_axi_mat_B_ch_1_AWADDR;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [1:0] m_axi_mat_B_ch_1_AWBURST;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [3:0] m_axi_mat_B_ch_1_AWCACHE;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [0:0] m_axi_mat_B_ch_1_AWID;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [7:0] m_axi_mat_B_ch_1_AWLEN;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output m_axi_mat_B_ch_1_AWLOCK;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [2:0] m_axi_mat_B_ch_1_AWPROT;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [3:0] m_axi_mat_B_ch_1_AWQOS;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.ready" *)input m_axi_mat_B_ch_1_AWREADY;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.data" *)output [2:0] m_axi_mat_B_ch_1_AWSIZE;
  (* RS_HS = "m_axi_mat_B_ch_1_AW.valid" *)output m_axi_mat_B_ch_1_AWVALID;
  (* RS_HS = "m_axi_mat_B_ch_1_B.data" *)input [0:0] m_axi_mat_B_ch_1_BID;
  (* RS_HS = "m_axi_mat_B_ch_1_B.ready" *)output m_axi_mat_B_ch_1_BREADY;
  (* RS_HS = "m_axi_mat_B_ch_1_B.data" *)input [1:0] m_axi_mat_B_ch_1_BRESP;
  (* RS_HS = "m_axi_mat_B_ch_1_B.valid" *)input m_axi_mat_B_ch_1_BVALID;
  (* RS_HS = "m_axi_mat_B_ch_1_R.data" *)input [511:0] m_axi_mat_B_ch_1_RDATA;
  (* RS_HS = "m_axi_mat_B_ch_1_R.data" *)input [0:0] m_axi_mat_B_ch_1_RID;
  (* RS_HS = "m_axi_mat_B_ch_1_R.data" *)input m_axi_mat_B_ch_1_RLAST;
  (* RS_HS = "m_axi_mat_B_ch_1_R.ready" *)output m_axi_mat_B_ch_1_RREADY;
  (* RS_HS = "m_axi_mat_B_ch_1_R.data" *)input [1:0] m_axi_mat_B_ch_1_RRESP;
  (* RS_HS = "m_axi_mat_B_ch_1_R.valid" *)input m_axi_mat_B_ch_1_RVALID;
  (* RS_HS = "m_axi_mat_B_ch_1_W.data" *)output [511:0] m_axi_mat_B_ch_1_WDATA;
  (* RS_HS = "m_axi_mat_B_ch_1_W.data" *)output m_axi_mat_B_ch_1_WLAST;
  (* RS_HS = "m_axi_mat_B_ch_1_W.ready" *)input m_axi_mat_B_ch_1_WREADY;
  (* RS_HS = "m_axi_mat_B_ch_1_W.data" *)output [63:0] m_axi_mat_B_ch_1_WSTRB;
  (* RS_HS = "m_axi_mat_B_ch_1_W.valid" *)output m_axi_mat_B_ch_1_WVALID;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [63:0] m_axi_mat_B_ch_2_ARADDR;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [1:0] m_axi_mat_B_ch_2_ARBURST;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [3:0] m_axi_mat_B_ch_2_ARCACHE;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [0:0] m_axi_mat_B_ch_2_ARID;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [7:0] m_axi_mat_B_ch_2_ARLEN;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output m_axi_mat_B_ch_2_ARLOCK;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [2:0] m_axi_mat_B_ch_2_ARPROT;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [3:0] m_axi_mat_B_ch_2_ARQOS;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.ready" *)input m_axi_mat_B_ch_2_ARREADY;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.data" *)output [2:0] m_axi_mat_B_ch_2_ARSIZE;
  (* RS_HS = "m_axi_mat_B_ch_2_AR.valid" *)output m_axi_mat_B_ch_2_ARVALID;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [63:0] m_axi_mat_B_ch_2_AWADDR;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [1:0] m_axi_mat_B_ch_2_AWBURST;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [3:0] m_axi_mat_B_ch_2_AWCACHE;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [0:0] m_axi_mat_B_ch_2_AWID;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [7:0] m_axi_mat_B_ch_2_AWLEN;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output m_axi_mat_B_ch_2_AWLOCK;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [2:0] m_axi_mat_B_ch_2_AWPROT;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [3:0] m_axi_mat_B_ch_2_AWQOS;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.ready" *)input m_axi_mat_B_ch_2_AWREADY;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.data" *)output [2:0] m_axi_mat_B_ch_2_AWSIZE;
  (* RS_HS = "m_axi_mat_B_ch_2_AW.valid" *)output m_axi_mat_B_ch_2_AWVALID;
  (* RS_HS = "m_axi_mat_B_ch_2_B.data" *)input [0:0] m_axi_mat_B_ch_2_BID;
  (* RS_HS = "m_axi_mat_B_ch_2_B.ready" *)output m_axi_mat_B_ch_2_BREADY;
  (* RS_HS = "m_axi_mat_B_ch_2_B.data" *)input [1:0] m_axi_mat_B_ch_2_BRESP;
  (* RS_HS = "m_axi_mat_B_ch_2_B.valid" *)input m_axi_mat_B_ch_2_BVALID;
  (* RS_HS = "m_axi_mat_B_ch_2_R.data" *)input [511:0] m_axi_mat_B_ch_2_RDATA;
  (* RS_HS = "m_axi_mat_B_ch_2_R.data" *)input [0:0] m_axi_mat_B_ch_2_RID;
  (* RS_HS = "m_axi_mat_B_ch_2_R.data" *)input m_axi_mat_B_ch_2_RLAST;
  (* RS_HS = "m_axi_mat_B_ch_2_R.ready" *)output m_axi_mat_B_ch_2_RREADY;
  (* RS_HS = "m_axi_mat_B_ch_2_R.data" *)input [1:0] m_axi_mat_B_ch_2_RRESP;
  (* RS_HS = "m_axi_mat_B_ch_2_R.valid" *)input m_axi_mat_B_ch_2_RVALID;
  (* RS_HS = "m_axi_mat_B_ch_2_W.data" *)output [511:0] m_axi_mat_B_ch_2_WDATA;
  (* RS_HS = "m_axi_mat_B_ch_2_W.data" *)output m_axi_mat_B_ch_2_WLAST;
  (* RS_HS = "m_axi_mat_B_ch_2_W.ready" *)input m_axi_mat_B_ch_2_WREADY;
  (* RS_HS = "m_axi_mat_B_ch_2_W.data" *)output [63:0] m_axi_mat_B_ch_2_WSTRB;
  (* RS_HS = "m_axi_mat_B_ch_2_W.valid" *)output m_axi_mat_B_ch_2_WVALID;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [63:0] m_axi_mat_B_ch_3_ARADDR;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [1:0] m_axi_mat_B_ch_3_ARBURST;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [3:0] m_axi_mat_B_ch_3_ARCACHE;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [0:0] m_axi_mat_B_ch_3_ARID;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [7:0] m_axi_mat_B_ch_3_ARLEN;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output m_axi_mat_B_ch_3_ARLOCK;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [2:0] m_axi_mat_B_ch_3_ARPROT;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [3:0] m_axi_mat_B_ch_3_ARQOS;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.ready" *)input m_axi_mat_B_ch_3_ARREADY;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.data" *)output [2:0] m_axi_mat_B_ch_3_ARSIZE;
  (* RS_HS = "m_axi_mat_B_ch_3_AR.valid" *)output m_axi_mat_B_ch_3_ARVALID;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [63:0] m_axi_mat_B_ch_3_AWADDR;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [1:0] m_axi_mat_B_ch_3_AWBURST;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [3:0] m_axi_mat_B_ch_3_AWCACHE;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [0:0] m_axi_mat_B_ch_3_AWID;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [7:0] m_axi_mat_B_ch_3_AWLEN;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output m_axi_mat_B_ch_3_AWLOCK;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [2:0] m_axi_mat_B_ch_3_AWPROT;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [3:0] m_axi_mat_B_ch_3_AWQOS;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.ready" *)input m_axi_mat_B_ch_3_AWREADY;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.data" *)output [2:0] m_axi_mat_B_ch_3_AWSIZE;
  (* RS_HS = "m_axi_mat_B_ch_3_AW.valid" *)output m_axi_mat_B_ch_3_AWVALID;
  (* RS_HS = "m_axi_mat_B_ch_3_B.data" *)input [0:0] m_axi_mat_B_ch_3_BID;
  (* RS_HS = "m_axi_mat_B_ch_3_B.ready" *)output m_axi_mat_B_ch_3_BREADY;
  (* RS_HS = "m_axi_mat_B_ch_3_B.data" *)input [1:0] m_axi_mat_B_ch_3_BRESP;
  (* RS_HS = "m_axi_mat_B_ch_3_B.valid" *)input m_axi_mat_B_ch_3_BVALID;
  (* RS_HS = "m_axi_mat_B_ch_3_R.data" *)input [511:0] m_axi_mat_B_ch_3_RDATA;
  (* RS_HS = "m_axi_mat_B_ch_3_R.data" *)input [0:0] m_axi_mat_B_ch_3_RID;
  (* RS_HS = "m_axi_mat_B_ch_3_R.data" *)input m_axi_mat_B_ch_3_RLAST;
  (* RS_HS = "m_axi_mat_B_ch_3_R.ready" *)output m_axi_mat_B_ch_3_RREADY;
  (* RS_HS = "m_axi_mat_B_ch_3_R.data" *)input [1:0] m_axi_mat_B_ch_3_RRESP;
  (* RS_HS = "m_axi_mat_B_ch_3_R.valid" *)input m_axi_mat_B_ch_3_RVALID;
  (* RS_HS = "m_axi_mat_B_ch_3_W.data" *)output [511:0] m_axi_mat_B_ch_3_WDATA;
  (* RS_HS = "m_axi_mat_B_ch_3_W.data" *)output m_axi_mat_B_ch_3_WLAST;
  (* RS_HS = "m_axi_mat_B_ch_3_W.ready" *)input m_axi_mat_B_ch_3_WREADY;
  (* RS_HS = "m_axi_mat_B_ch_3_W.data" *)output [63:0] m_axi_mat_B_ch_3_WSTRB;
  (* RS_HS = "m_axi_mat_B_ch_3_W.valid" *)output m_axi_mat_B_ch_3_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [63:0] m_axi_mat_C_ch_in_0_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [1:0] m_axi_mat_C_ch_in_0_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [3:0] m_axi_mat_C_ch_in_0_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [0:0] m_axi_mat_C_ch_in_0_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [7:0] m_axi_mat_C_ch_in_0_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output m_axi_mat_C_ch_in_0_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [2:0] m_axi_mat_C_ch_in_0_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [3:0] m_axi_mat_C_ch_in_0_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.ready" *)input m_axi_mat_C_ch_in_0_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.data" *)output [2:0] m_axi_mat_C_ch_in_0_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AR.valid" *)output m_axi_mat_C_ch_in_0_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [63:0] m_axi_mat_C_ch_in_0_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [1:0] m_axi_mat_C_ch_in_0_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [3:0] m_axi_mat_C_ch_in_0_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [0:0] m_axi_mat_C_ch_in_0_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [7:0] m_axi_mat_C_ch_in_0_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output m_axi_mat_C_ch_in_0_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [2:0] m_axi_mat_C_ch_in_0_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [3:0] m_axi_mat_C_ch_in_0_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.ready" *)input m_axi_mat_C_ch_in_0_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.data" *)output [2:0] m_axi_mat_C_ch_in_0_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_0_AW.valid" *)output m_axi_mat_C_ch_in_0_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_B.data" *)input [0:0] m_axi_mat_C_ch_in_0_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_B.ready" *)output m_axi_mat_C_ch_in_0_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_0_B.data" *)input [1:0] m_axi_mat_C_ch_in_0_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_0_B.valid" *)input m_axi_mat_C_ch_in_0_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_R.data" *)input [511:0] m_axi_mat_C_ch_in_0_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_0_R.data" *)input [0:0] m_axi_mat_C_ch_in_0_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_R.data" *)input m_axi_mat_C_ch_in_0_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_0_R.ready" *)output m_axi_mat_C_ch_in_0_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_0_R.data" *)input [1:0] m_axi_mat_C_ch_in_0_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_0_R.valid" *)input m_axi_mat_C_ch_in_0_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_0_W.data" *)output [511:0] m_axi_mat_C_ch_in_0_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_0_W.data" *)output m_axi_mat_C_ch_in_0_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_0_W.ready" *)input m_axi_mat_C_ch_in_0_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_0_W.data" *)output [63:0] m_axi_mat_C_ch_in_0_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_0_W.valid" *)output m_axi_mat_C_ch_in_0_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [63:0] m_axi_mat_C_ch_in_1_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [1:0] m_axi_mat_C_ch_in_1_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [3:0] m_axi_mat_C_ch_in_1_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [0:0] m_axi_mat_C_ch_in_1_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [7:0] m_axi_mat_C_ch_in_1_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output m_axi_mat_C_ch_in_1_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [2:0] m_axi_mat_C_ch_in_1_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [3:0] m_axi_mat_C_ch_in_1_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.ready" *)input m_axi_mat_C_ch_in_1_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.data" *)output [2:0] m_axi_mat_C_ch_in_1_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AR.valid" *)output m_axi_mat_C_ch_in_1_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [63:0] m_axi_mat_C_ch_in_1_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [1:0] m_axi_mat_C_ch_in_1_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [3:0] m_axi_mat_C_ch_in_1_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [0:0] m_axi_mat_C_ch_in_1_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [7:0] m_axi_mat_C_ch_in_1_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output m_axi_mat_C_ch_in_1_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [2:0] m_axi_mat_C_ch_in_1_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [3:0] m_axi_mat_C_ch_in_1_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.ready" *)input m_axi_mat_C_ch_in_1_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.data" *)output [2:0] m_axi_mat_C_ch_in_1_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_1_AW.valid" *)output m_axi_mat_C_ch_in_1_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_B.data" *)input [0:0] m_axi_mat_C_ch_in_1_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_B.ready" *)output m_axi_mat_C_ch_in_1_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_1_B.data" *)input [1:0] m_axi_mat_C_ch_in_1_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_1_B.valid" *)input m_axi_mat_C_ch_in_1_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_R.data" *)input [511:0] m_axi_mat_C_ch_in_1_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_1_R.data" *)input [0:0] m_axi_mat_C_ch_in_1_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_R.data" *)input m_axi_mat_C_ch_in_1_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_1_R.ready" *)output m_axi_mat_C_ch_in_1_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_1_R.data" *)input [1:0] m_axi_mat_C_ch_in_1_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_1_R.valid" *)input m_axi_mat_C_ch_in_1_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_1_W.data" *)output [511:0] m_axi_mat_C_ch_in_1_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_1_W.data" *)output m_axi_mat_C_ch_in_1_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_1_W.ready" *)input m_axi_mat_C_ch_in_1_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_1_W.data" *)output [63:0] m_axi_mat_C_ch_in_1_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_1_W.valid" *)output m_axi_mat_C_ch_in_1_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [63:0] m_axi_mat_C_ch_in_2_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [1:0] m_axi_mat_C_ch_in_2_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [3:0] m_axi_mat_C_ch_in_2_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [0:0] m_axi_mat_C_ch_in_2_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [7:0] m_axi_mat_C_ch_in_2_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output m_axi_mat_C_ch_in_2_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [2:0] m_axi_mat_C_ch_in_2_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [3:0] m_axi_mat_C_ch_in_2_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.ready" *)input m_axi_mat_C_ch_in_2_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.data" *)output [2:0] m_axi_mat_C_ch_in_2_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AR.valid" *)output m_axi_mat_C_ch_in_2_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [63:0] m_axi_mat_C_ch_in_2_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [1:0] m_axi_mat_C_ch_in_2_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [3:0] m_axi_mat_C_ch_in_2_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [0:0] m_axi_mat_C_ch_in_2_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [7:0] m_axi_mat_C_ch_in_2_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output m_axi_mat_C_ch_in_2_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [2:0] m_axi_mat_C_ch_in_2_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [3:0] m_axi_mat_C_ch_in_2_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.ready" *)input m_axi_mat_C_ch_in_2_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.data" *)output [2:0] m_axi_mat_C_ch_in_2_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_2_AW.valid" *)output m_axi_mat_C_ch_in_2_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_B.data" *)input [0:0] m_axi_mat_C_ch_in_2_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_B.ready" *)output m_axi_mat_C_ch_in_2_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_2_B.data" *)input [1:0] m_axi_mat_C_ch_in_2_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_2_B.valid" *)input m_axi_mat_C_ch_in_2_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_R.data" *)input [511:0] m_axi_mat_C_ch_in_2_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_2_R.data" *)input [0:0] m_axi_mat_C_ch_in_2_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_R.data" *)input m_axi_mat_C_ch_in_2_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_2_R.ready" *)output m_axi_mat_C_ch_in_2_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_2_R.data" *)input [1:0] m_axi_mat_C_ch_in_2_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_2_R.valid" *)input m_axi_mat_C_ch_in_2_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_2_W.data" *)output [511:0] m_axi_mat_C_ch_in_2_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_2_W.data" *)output m_axi_mat_C_ch_in_2_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_2_W.ready" *)input m_axi_mat_C_ch_in_2_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_2_W.data" *)output [63:0] m_axi_mat_C_ch_in_2_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_2_W.valid" *)output m_axi_mat_C_ch_in_2_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [63:0] m_axi_mat_C_ch_in_3_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [1:0] m_axi_mat_C_ch_in_3_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [3:0] m_axi_mat_C_ch_in_3_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [0:0] m_axi_mat_C_ch_in_3_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [7:0] m_axi_mat_C_ch_in_3_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output m_axi_mat_C_ch_in_3_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [2:0] m_axi_mat_C_ch_in_3_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [3:0] m_axi_mat_C_ch_in_3_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.ready" *)input m_axi_mat_C_ch_in_3_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.data" *)output [2:0] m_axi_mat_C_ch_in_3_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AR.valid" *)output m_axi_mat_C_ch_in_3_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [63:0] m_axi_mat_C_ch_in_3_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [1:0] m_axi_mat_C_ch_in_3_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [3:0] m_axi_mat_C_ch_in_3_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [0:0] m_axi_mat_C_ch_in_3_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [7:0] m_axi_mat_C_ch_in_3_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output m_axi_mat_C_ch_in_3_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [2:0] m_axi_mat_C_ch_in_3_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [3:0] m_axi_mat_C_ch_in_3_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.ready" *)input m_axi_mat_C_ch_in_3_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.data" *)output [2:0] m_axi_mat_C_ch_in_3_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_3_AW.valid" *)output m_axi_mat_C_ch_in_3_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_B.data" *)input [0:0] m_axi_mat_C_ch_in_3_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_B.ready" *)output m_axi_mat_C_ch_in_3_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_3_B.data" *)input [1:0] m_axi_mat_C_ch_in_3_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_3_B.valid" *)input m_axi_mat_C_ch_in_3_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_R.data" *)input [511:0] m_axi_mat_C_ch_in_3_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_3_R.data" *)input [0:0] m_axi_mat_C_ch_in_3_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_R.data" *)input m_axi_mat_C_ch_in_3_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_3_R.ready" *)output m_axi_mat_C_ch_in_3_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_3_R.data" *)input [1:0] m_axi_mat_C_ch_in_3_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_3_R.valid" *)input m_axi_mat_C_ch_in_3_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_3_W.data" *)output [511:0] m_axi_mat_C_ch_in_3_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_3_W.data" *)output m_axi_mat_C_ch_in_3_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_3_W.ready" *)input m_axi_mat_C_ch_in_3_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_3_W.data" *)output [63:0] m_axi_mat_C_ch_in_3_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_3_W.valid" *)output m_axi_mat_C_ch_in_3_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [63:0] m_axi_mat_C_ch_in_4_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [1:0] m_axi_mat_C_ch_in_4_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [3:0] m_axi_mat_C_ch_in_4_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [0:0] m_axi_mat_C_ch_in_4_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [7:0] m_axi_mat_C_ch_in_4_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output m_axi_mat_C_ch_in_4_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [2:0] m_axi_mat_C_ch_in_4_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [3:0] m_axi_mat_C_ch_in_4_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.ready" *)input m_axi_mat_C_ch_in_4_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.data" *)output [2:0] m_axi_mat_C_ch_in_4_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AR.valid" *)output m_axi_mat_C_ch_in_4_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [63:0] m_axi_mat_C_ch_in_4_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [1:0] m_axi_mat_C_ch_in_4_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [3:0] m_axi_mat_C_ch_in_4_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [0:0] m_axi_mat_C_ch_in_4_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [7:0] m_axi_mat_C_ch_in_4_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output m_axi_mat_C_ch_in_4_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [2:0] m_axi_mat_C_ch_in_4_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [3:0] m_axi_mat_C_ch_in_4_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.ready" *)input m_axi_mat_C_ch_in_4_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.data" *)output [2:0] m_axi_mat_C_ch_in_4_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_4_AW.valid" *)output m_axi_mat_C_ch_in_4_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_B.data" *)input [0:0] m_axi_mat_C_ch_in_4_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_B.ready" *)output m_axi_mat_C_ch_in_4_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_4_B.data" *)input [1:0] m_axi_mat_C_ch_in_4_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_4_B.valid" *)input m_axi_mat_C_ch_in_4_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_R.data" *)input [511:0] m_axi_mat_C_ch_in_4_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_4_R.data" *)input [0:0] m_axi_mat_C_ch_in_4_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_R.data" *)input m_axi_mat_C_ch_in_4_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_4_R.ready" *)output m_axi_mat_C_ch_in_4_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_4_R.data" *)input [1:0] m_axi_mat_C_ch_in_4_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_4_R.valid" *)input m_axi_mat_C_ch_in_4_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_4_W.data" *)output [511:0] m_axi_mat_C_ch_in_4_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_4_W.data" *)output m_axi_mat_C_ch_in_4_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_4_W.ready" *)input m_axi_mat_C_ch_in_4_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_4_W.data" *)output [63:0] m_axi_mat_C_ch_in_4_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_4_W.valid" *)output m_axi_mat_C_ch_in_4_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [63:0] m_axi_mat_C_ch_in_5_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [1:0] m_axi_mat_C_ch_in_5_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [3:0] m_axi_mat_C_ch_in_5_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [0:0] m_axi_mat_C_ch_in_5_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [7:0] m_axi_mat_C_ch_in_5_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output m_axi_mat_C_ch_in_5_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [2:0] m_axi_mat_C_ch_in_5_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [3:0] m_axi_mat_C_ch_in_5_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.ready" *)input m_axi_mat_C_ch_in_5_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.data" *)output [2:0] m_axi_mat_C_ch_in_5_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AR.valid" *)output m_axi_mat_C_ch_in_5_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [63:0] m_axi_mat_C_ch_in_5_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [1:0] m_axi_mat_C_ch_in_5_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [3:0] m_axi_mat_C_ch_in_5_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [0:0] m_axi_mat_C_ch_in_5_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [7:0] m_axi_mat_C_ch_in_5_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output m_axi_mat_C_ch_in_5_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [2:0] m_axi_mat_C_ch_in_5_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [3:0] m_axi_mat_C_ch_in_5_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.ready" *)input m_axi_mat_C_ch_in_5_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.data" *)output [2:0] m_axi_mat_C_ch_in_5_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_5_AW.valid" *)output m_axi_mat_C_ch_in_5_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_B.data" *)input [0:0] m_axi_mat_C_ch_in_5_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_B.ready" *)output m_axi_mat_C_ch_in_5_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_5_B.data" *)input [1:0] m_axi_mat_C_ch_in_5_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_5_B.valid" *)input m_axi_mat_C_ch_in_5_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_R.data" *)input [511:0] m_axi_mat_C_ch_in_5_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_5_R.data" *)input [0:0] m_axi_mat_C_ch_in_5_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_R.data" *)input m_axi_mat_C_ch_in_5_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_5_R.ready" *)output m_axi_mat_C_ch_in_5_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_5_R.data" *)input [1:0] m_axi_mat_C_ch_in_5_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_5_R.valid" *)input m_axi_mat_C_ch_in_5_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_5_W.data" *)output [511:0] m_axi_mat_C_ch_in_5_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_5_W.data" *)output m_axi_mat_C_ch_in_5_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_5_W.ready" *)input m_axi_mat_C_ch_in_5_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_5_W.data" *)output [63:0] m_axi_mat_C_ch_in_5_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_5_W.valid" *)output m_axi_mat_C_ch_in_5_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [63:0] m_axi_mat_C_ch_in_6_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [1:0] m_axi_mat_C_ch_in_6_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [3:0] m_axi_mat_C_ch_in_6_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [0:0] m_axi_mat_C_ch_in_6_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [7:0] m_axi_mat_C_ch_in_6_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output m_axi_mat_C_ch_in_6_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [2:0] m_axi_mat_C_ch_in_6_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [3:0] m_axi_mat_C_ch_in_6_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.ready" *)input m_axi_mat_C_ch_in_6_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.data" *)output [2:0] m_axi_mat_C_ch_in_6_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AR.valid" *)output m_axi_mat_C_ch_in_6_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [63:0] m_axi_mat_C_ch_in_6_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [1:0] m_axi_mat_C_ch_in_6_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [3:0] m_axi_mat_C_ch_in_6_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [0:0] m_axi_mat_C_ch_in_6_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [7:0] m_axi_mat_C_ch_in_6_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output m_axi_mat_C_ch_in_6_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [2:0] m_axi_mat_C_ch_in_6_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [3:0] m_axi_mat_C_ch_in_6_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.ready" *)input m_axi_mat_C_ch_in_6_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.data" *)output [2:0] m_axi_mat_C_ch_in_6_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_6_AW.valid" *)output m_axi_mat_C_ch_in_6_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_B.data" *)input [0:0] m_axi_mat_C_ch_in_6_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_B.ready" *)output m_axi_mat_C_ch_in_6_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_6_B.data" *)input [1:0] m_axi_mat_C_ch_in_6_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_6_B.valid" *)input m_axi_mat_C_ch_in_6_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_R.data" *)input [511:0] m_axi_mat_C_ch_in_6_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_6_R.data" *)input [0:0] m_axi_mat_C_ch_in_6_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_R.data" *)input m_axi_mat_C_ch_in_6_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_6_R.ready" *)output m_axi_mat_C_ch_in_6_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_6_R.data" *)input [1:0] m_axi_mat_C_ch_in_6_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_6_R.valid" *)input m_axi_mat_C_ch_in_6_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_6_W.data" *)output [511:0] m_axi_mat_C_ch_in_6_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_6_W.data" *)output m_axi_mat_C_ch_in_6_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_6_W.ready" *)input m_axi_mat_C_ch_in_6_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_6_W.data" *)output [63:0] m_axi_mat_C_ch_in_6_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_6_W.valid" *)output m_axi_mat_C_ch_in_6_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [63:0] m_axi_mat_C_ch_in_7_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [1:0] m_axi_mat_C_ch_in_7_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [3:0] m_axi_mat_C_ch_in_7_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [0:0] m_axi_mat_C_ch_in_7_ARID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [7:0] m_axi_mat_C_ch_in_7_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output m_axi_mat_C_ch_in_7_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [2:0] m_axi_mat_C_ch_in_7_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [3:0] m_axi_mat_C_ch_in_7_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.ready" *)input m_axi_mat_C_ch_in_7_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.data" *)output [2:0] m_axi_mat_C_ch_in_7_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AR.valid" *)output m_axi_mat_C_ch_in_7_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [63:0] m_axi_mat_C_ch_in_7_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [1:0] m_axi_mat_C_ch_in_7_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [3:0] m_axi_mat_C_ch_in_7_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [0:0] m_axi_mat_C_ch_in_7_AWID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [7:0] m_axi_mat_C_ch_in_7_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output m_axi_mat_C_ch_in_7_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [2:0] m_axi_mat_C_ch_in_7_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [3:0] m_axi_mat_C_ch_in_7_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.ready" *)input m_axi_mat_C_ch_in_7_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.data" *)output [2:0] m_axi_mat_C_ch_in_7_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_in_7_AW.valid" *)output m_axi_mat_C_ch_in_7_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_B.data" *)input [0:0] m_axi_mat_C_ch_in_7_BID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_B.ready" *)output m_axi_mat_C_ch_in_7_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_7_B.data" *)input [1:0] m_axi_mat_C_ch_in_7_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_7_B.valid" *)input m_axi_mat_C_ch_in_7_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_R.data" *)input [511:0] m_axi_mat_C_ch_in_7_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_7_R.data" *)input [0:0] m_axi_mat_C_ch_in_7_RID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_R.data" *)input m_axi_mat_C_ch_in_7_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_7_R.ready" *)output m_axi_mat_C_ch_in_7_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_7_R.data" *)input [1:0] m_axi_mat_C_ch_in_7_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_in_7_R.valid" *)input m_axi_mat_C_ch_in_7_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_in_7_W.data" *)output [511:0] m_axi_mat_C_ch_in_7_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_in_7_W.data" *)output m_axi_mat_C_ch_in_7_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_in_7_W.ready" *)input m_axi_mat_C_ch_in_7_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_in_7_W.data" *)output [63:0] m_axi_mat_C_ch_in_7_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_in_7_W.valid" *)output m_axi_mat_C_ch_in_7_WVALID;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [63:0] m_axi_edge_list_ptr_ARADDR;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [1:0] m_axi_edge_list_ptr_ARBURST;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [3:0] m_axi_edge_list_ptr_ARCACHE;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [0:0] m_axi_edge_list_ptr_ARID;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [7:0] m_axi_edge_list_ptr_ARLEN;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output m_axi_edge_list_ptr_ARLOCK;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [2:0] m_axi_edge_list_ptr_ARPROT;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [3:0] m_axi_edge_list_ptr_ARQOS;
  (* RS_HS = "m_axi_edge_list_ptr_AR.ready" *)input m_axi_edge_list_ptr_ARREADY;
  (* RS_HS = "m_axi_edge_list_ptr_AR.data" *)output [2:0] m_axi_edge_list_ptr_ARSIZE;
  (* RS_HS = "m_axi_edge_list_ptr_AR.valid" *)output m_axi_edge_list_ptr_ARVALID;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [63:0] m_axi_edge_list_ptr_AWADDR;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [1:0] m_axi_edge_list_ptr_AWBURST;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [3:0] m_axi_edge_list_ptr_AWCACHE;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [0:0] m_axi_edge_list_ptr_AWID;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [7:0] m_axi_edge_list_ptr_AWLEN;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output m_axi_edge_list_ptr_AWLOCK;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [2:0] m_axi_edge_list_ptr_AWPROT;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [3:0] m_axi_edge_list_ptr_AWQOS;
  (* RS_HS = "m_axi_edge_list_ptr_AW.ready" *)input m_axi_edge_list_ptr_AWREADY;
  (* RS_HS = "m_axi_edge_list_ptr_AW.data" *)output [2:0] m_axi_edge_list_ptr_AWSIZE;
  (* RS_HS = "m_axi_edge_list_ptr_AW.valid" *)output m_axi_edge_list_ptr_AWVALID;
  (* RS_HS = "m_axi_edge_list_ptr_B.data" *)input [0:0] m_axi_edge_list_ptr_BID;
  (* RS_HS = "m_axi_edge_list_ptr_B.ready" *)output m_axi_edge_list_ptr_BREADY;
  (* RS_HS = "m_axi_edge_list_ptr_B.data" *)input [1:0] m_axi_edge_list_ptr_BRESP;
  (* RS_HS = "m_axi_edge_list_ptr_B.valid" *)input m_axi_edge_list_ptr_BVALID;
  (* RS_HS = "m_axi_edge_list_ptr_R.data" *)input [31:0] m_axi_edge_list_ptr_RDATA;
  (* RS_HS = "m_axi_edge_list_ptr_R.data" *)input [0:0] m_axi_edge_list_ptr_RID;
  (* RS_HS = "m_axi_edge_list_ptr_R.data" *)input m_axi_edge_list_ptr_RLAST;
  (* RS_HS = "m_axi_edge_list_ptr_R.ready" *)output m_axi_edge_list_ptr_RREADY;
  (* RS_HS = "m_axi_edge_list_ptr_R.data" *)input [1:0] m_axi_edge_list_ptr_RRESP;
  (* RS_HS = "m_axi_edge_list_ptr_R.valid" *)input m_axi_edge_list_ptr_RVALID;
  (* RS_HS = "m_axi_edge_list_ptr_W.data" *)output [31:0] m_axi_edge_list_ptr_WDATA;
  (* RS_HS = "m_axi_edge_list_ptr_W.data" *)output m_axi_edge_list_ptr_WLAST;
  (* RS_HS = "m_axi_edge_list_ptr_W.ready" *)input m_axi_edge_list_ptr_WREADY;
  (* RS_HS = "m_axi_edge_list_ptr_W.data" *)output [3:0] m_axi_edge_list_ptr_WSTRB;
  (* RS_HS = "m_axi_edge_list_ptr_W.valid" *)output m_axi_edge_list_ptr_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [63:0] m_axi_mat_C_ch_0_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [1:0] m_axi_mat_C_ch_0_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [3:0] m_axi_mat_C_ch_0_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [0:0] m_axi_mat_C_ch_0_ARID;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [7:0] m_axi_mat_C_ch_0_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output m_axi_mat_C_ch_0_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [2:0] m_axi_mat_C_ch_0_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [3:0] m_axi_mat_C_ch_0_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.ready" *)input m_axi_mat_C_ch_0_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.data" *)output [2:0] m_axi_mat_C_ch_0_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_0_AR.valid" *)output m_axi_mat_C_ch_0_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [63:0] m_axi_mat_C_ch_0_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [1:0] m_axi_mat_C_ch_0_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [3:0] m_axi_mat_C_ch_0_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [0:0] m_axi_mat_C_ch_0_AWID;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [7:0] m_axi_mat_C_ch_0_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output m_axi_mat_C_ch_0_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [2:0] m_axi_mat_C_ch_0_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [3:0] m_axi_mat_C_ch_0_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.ready" *)input m_axi_mat_C_ch_0_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.data" *)output [2:0] m_axi_mat_C_ch_0_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_0_AW.valid" *)output m_axi_mat_C_ch_0_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_0_B.data" *)input [0:0] m_axi_mat_C_ch_0_BID;
  (* RS_HS = "m_axi_mat_C_ch_0_B.ready" *)output m_axi_mat_C_ch_0_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_0_B.data" *)input [1:0] m_axi_mat_C_ch_0_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_0_B.valid" *)input m_axi_mat_C_ch_0_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_0_R.data" *)input [511:0] m_axi_mat_C_ch_0_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_0_R.data" *)input [0:0] m_axi_mat_C_ch_0_RID;
  (* RS_HS = "m_axi_mat_C_ch_0_R.data" *)input m_axi_mat_C_ch_0_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_0_R.ready" *)output m_axi_mat_C_ch_0_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_0_R.data" *)input [1:0] m_axi_mat_C_ch_0_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_0_R.valid" *)input m_axi_mat_C_ch_0_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_0_W.data" *)output [511:0] m_axi_mat_C_ch_0_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_0_W.data" *)output m_axi_mat_C_ch_0_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_0_W.ready" *)input m_axi_mat_C_ch_0_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_0_W.data" *)output [63:0] m_axi_mat_C_ch_0_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_0_W.valid" *)output m_axi_mat_C_ch_0_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [63:0] m_axi_mat_C_ch_1_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [1:0] m_axi_mat_C_ch_1_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [3:0] m_axi_mat_C_ch_1_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [0:0] m_axi_mat_C_ch_1_ARID;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [7:0] m_axi_mat_C_ch_1_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output m_axi_mat_C_ch_1_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [2:0] m_axi_mat_C_ch_1_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [3:0] m_axi_mat_C_ch_1_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.ready" *)input m_axi_mat_C_ch_1_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.data" *)output [2:0] m_axi_mat_C_ch_1_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_1_AR.valid" *)output m_axi_mat_C_ch_1_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [63:0] m_axi_mat_C_ch_1_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [1:0] m_axi_mat_C_ch_1_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [3:0] m_axi_mat_C_ch_1_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [0:0] m_axi_mat_C_ch_1_AWID;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [7:0] m_axi_mat_C_ch_1_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output m_axi_mat_C_ch_1_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [2:0] m_axi_mat_C_ch_1_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [3:0] m_axi_mat_C_ch_1_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.ready" *)input m_axi_mat_C_ch_1_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.data" *)output [2:0] m_axi_mat_C_ch_1_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_1_AW.valid" *)output m_axi_mat_C_ch_1_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_1_B.data" *)input [0:0] m_axi_mat_C_ch_1_BID;
  (* RS_HS = "m_axi_mat_C_ch_1_B.ready" *)output m_axi_mat_C_ch_1_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_1_B.data" *)input [1:0] m_axi_mat_C_ch_1_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_1_B.valid" *)input m_axi_mat_C_ch_1_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_1_R.data" *)input [511:0] m_axi_mat_C_ch_1_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_1_R.data" *)input [0:0] m_axi_mat_C_ch_1_RID;
  (* RS_HS = "m_axi_mat_C_ch_1_R.data" *)input m_axi_mat_C_ch_1_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_1_R.ready" *)output m_axi_mat_C_ch_1_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_1_R.data" *)input [1:0] m_axi_mat_C_ch_1_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_1_R.valid" *)input m_axi_mat_C_ch_1_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_1_W.data" *)output [511:0] m_axi_mat_C_ch_1_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_1_W.data" *)output m_axi_mat_C_ch_1_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_1_W.ready" *)input m_axi_mat_C_ch_1_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_1_W.data" *)output [63:0] m_axi_mat_C_ch_1_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_1_W.valid" *)output m_axi_mat_C_ch_1_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [63:0] m_axi_mat_C_ch_2_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [1:0] m_axi_mat_C_ch_2_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [3:0] m_axi_mat_C_ch_2_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [0:0] m_axi_mat_C_ch_2_ARID;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [7:0] m_axi_mat_C_ch_2_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output m_axi_mat_C_ch_2_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [2:0] m_axi_mat_C_ch_2_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [3:0] m_axi_mat_C_ch_2_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.ready" *)input m_axi_mat_C_ch_2_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.data" *)output [2:0] m_axi_mat_C_ch_2_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_2_AR.valid" *)output m_axi_mat_C_ch_2_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [63:0] m_axi_mat_C_ch_2_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [1:0] m_axi_mat_C_ch_2_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [3:0] m_axi_mat_C_ch_2_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [0:0] m_axi_mat_C_ch_2_AWID;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [7:0] m_axi_mat_C_ch_2_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output m_axi_mat_C_ch_2_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [2:0] m_axi_mat_C_ch_2_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [3:0] m_axi_mat_C_ch_2_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.ready" *)input m_axi_mat_C_ch_2_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.data" *)output [2:0] m_axi_mat_C_ch_2_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_2_AW.valid" *)output m_axi_mat_C_ch_2_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_2_B.data" *)input [0:0] m_axi_mat_C_ch_2_BID;
  (* RS_HS = "m_axi_mat_C_ch_2_B.ready" *)output m_axi_mat_C_ch_2_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_2_B.data" *)input [1:0] m_axi_mat_C_ch_2_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_2_B.valid" *)input m_axi_mat_C_ch_2_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_2_R.data" *)input [511:0] m_axi_mat_C_ch_2_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_2_R.data" *)input [0:0] m_axi_mat_C_ch_2_RID;
  (* RS_HS = "m_axi_mat_C_ch_2_R.data" *)input m_axi_mat_C_ch_2_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_2_R.ready" *)output m_axi_mat_C_ch_2_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_2_R.data" *)input [1:0] m_axi_mat_C_ch_2_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_2_R.valid" *)input m_axi_mat_C_ch_2_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_2_W.data" *)output [511:0] m_axi_mat_C_ch_2_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_2_W.data" *)output m_axi_mat_C_ch_2_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_2_W.ready" *)input m_axi_mat_C_ch_2_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_2_W.data" *)output [63:0] m_axi_mat_C_ch_2_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_2_W.valid" *)output m_axi_mat_C_ch_2_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [63:0] m_axi_mat_C_ch_3_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [1:0] m_axi_mat_C_ch_3_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [3:0] m_axi_mat_C_ch_3_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [0:0] m_axi_mat_C_ch_3_ARID;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [7:0] m_axi_mat_C_ch_3_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output m_axi_mat_C_ch_3_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [2:0] m_axi_mat_C_ch_3_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [3:0] m_axi_mat_C_ch_3_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.ready" *)input m_axi_mat_C_ch_3_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.data" *)output [2:0] m_axi_mat_C_ch_3_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_3_AR.valid" *)output m_axi_mat_C_ch_3_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [63:0] m_axi_mat_C_ch_3_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [1:0] m_axi_mat_C_ch_3_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [3:0] m_axi_mat_C_ch_3_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [0:0] m_axi_mat_C_ch_3_AWID;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [7:0] m_axi_mat_C_ch_3_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output m_axi_mat_C_ch_3_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [2:0] m_axi_mat_C_ch_3_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [3:0] m_axi_mat_C_ch_3_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.ready" *)input m_axi_mat_C_ch_3_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.data" *)output [2:0] m_axi_mat_C_ch_3_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_3_AW.valid" *)output m_axi_mat_C_ch_3_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_3_B.data" *)input [0:0] m_axi_mat_C_ch_3_BID;
  (* RS_HS = "m_axi_mat_C_ch_3_B.ready" *)output m_axi_mat_C_ch_3_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_3_B.data" *)input [1:0] m_axi_mat_C_ch_3_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_3_B.valid" *)input m_axi_mat_C_ch_3_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_3_R.data" *)input [511:0] m_axi_mat_C_ch_3_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_3_R.data" *)input [0:0] m_axi_mat_C_ch_3_RID;
  (* RS_HS = "m_axi_mat_C_ch_3_R.data" *)input m_axi_mat_C_ch_3_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_3_R.ready" *)output m_axi_mat_C_ch_3_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_3_R.data" *)input [1:0] m_axi_mat_C_ch_3_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_3_R.valid" *)input m_axi_mat_C_ch_3_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_3_W.data" *)output [511:0] m_axi_mat_C_ch_3_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_3_W.data" *)output m_axi_mat_C_ch_3_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_3_W.ready" *)input m_axi_mat_C_ch_3_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_3_W.data" *)output [63:0] m_axi_mat_C_ch_3_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_3_W.valid" *)output m_axi_mat_C_ch_3_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [63:0] m_axi_mat_C_ch_4_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [1:0] m_axi_mat_C_ch_4_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [3:0] m_axi_mat_C_ch_4_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [0:0] m_axi_mat_C_ch_4_ARID;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [7:0] m_axi_mat_C_ch_4_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output m_axi_mat_C_ch_4_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [2:0] m_axi_mat_C_ch_4_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [3:0] m_axi_mat_C_ch_4_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.ready" *)input m_axi_mat_C_ch_4_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.data" *)output [2:0] m_axi_mat_C_ch_4_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_4_AR.valid" *)output m_axi_mat_C_ch_4_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [63:0] m_axi_mat_C_ch_4_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [1:0] m_axi_mat_C_ch_4_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [3:0] m_axi_mat_C_ch_4_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [0:0] m_axi_mat_C_ch_4_AWID;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [7:0] m_axi_mat_C_ch_4_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output m_axi_mat_C_ch_4_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [2:0] m_axi_mat_C_ch_4_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [3:0] m_axi_mat_C_ch_4_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.ready" *)input m_axi_mat_C_ch_4_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.data" *)output [2:0] m_axi_mat_C_ch_4_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_4_AW.valid" *)output m_axi_mat_C_ch_4_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_4_B.data" *)input [0:0] m_axi_mat_C_ch_4_BID;
  (* RS_HS = "m_axi_mat_C_ch_4_B.ready" *)output m_axi_mat_C_ch_4_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_4_B.data" *)input [1:0] m_axi_mat_C_ch_4_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_4_B.valid" *)input m_axi_mat_C_ch_4_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_4_R.data" *)input [511:0] m_axi_mat_C_ch_4_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_4_R.data" *)input [0:0] m_axi_mat_C_ch_4_RID;
  (* RS_HS = "m_axi_mat_C_ch_4_R.data" *)input m_axi_mat_C_ch_4_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_4_R.ready" *)output m_axi_mat_C_ch_4_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_4_R.data" *)input [1:0] m_axi_mat_C_ch_4_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_4_R.valid" *)input m_axi_mat_C_ch_4_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_4_W.data" *)output [511:0] m_axi_mat_C_ch_4_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_4_W.data" *)output m_axi_mat_C_ch_4_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_4_W.ready" *)input m_axi_mat_C_ch_4_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_4_W.data" *)output [63:0] m_axi_mat_C_ch_4_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_4_W.valid" *)output m_axi_mat_C_ch_4_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [63:0] m_axi_mat_C_ch_5_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [1:0] m_axi_mat_C_ch_5_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [3:0] m_axi_mat_C_ch_5_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [0:0] m_axi_mat_C_ch_5_ARID;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [7:0] m_axi_mat_C_ch_5_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output m_axi_mat_C_ch_5_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [2:0] m_axi_mat_C_ch_5_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [3:0] m_axi_mat_C_ch_5_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.ready" *)input m_axi_mat_C_ch_5_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.data" *)output [2:0] m_axi_mat_C_ch_5_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_5_AR.valid" *)output m_axi_mat_C_ch_5_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [63:0] m_axi_mat_C_ch_5_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [1:0] m_axi_mat_C_ch_5_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [3:0] m_axi_mat_C_ch_5_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [0:0] m_axi_mat_C_ch_5_AWID;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [7:0] m_axi_mat_C_ch_5_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output m_axi_mat_C_ch_5_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [2:0] m_axi_mat_C_ch_5_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [3:0] m_axi_mat_C_ch_5_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.ready" *)input m_axi_mat_C_ch_5_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.data" *)output [2:0] m_axi_mat_C_ch_5_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_5_AW.valid" *)output m_axi_mat_C_ch_5_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_5_B.data" *)input [0:0] m_axi_mat_C_ch_5_BID;
  (* RS_HS = "m_axi_mat_C_ch_5_B.ready" *)output m_axi_mat_C_ch_5_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_5_B.data" *)input [1:0] m_axi_mat_C_ch_5_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_5_B.valid" *)input m_axi_mat_C_ch_5_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_5_R.data" *)input [511:0] m_axi_mat_C_ch_5_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_5_R.data" *)input [0:0] m_axi_mat_C_ch_5_RID;
  (* RS_HS = "m_axi_mat_C_ch_5_R.data" *)input m_axi_mat_C_ch_5_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_5_R.ready" *)output m_axi_mat_C_ch_5_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_5_R.data" *)input [1:0] m_axi_mat_C_ch_5_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_5_R.valid" *)input m_axi_mat_C_ch_5_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_5_W.data" *)output [511:0] m_axi_mat_C_ch_5_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_5_W.data" *)output m_axi_mat_C_ch_5_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_5_W.ready" *)input m_axi_mat_C_ch_5_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_5_W.data" *)output [63:0] m_axi_mat_C_ch_5_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_5_W.valid" *)output m_axi_mat_C_ch_5_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [63:0] m_axi_mat_C_ch_6_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [1:0] m_axi_mat_C_ch_6_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [3:0] m_axi_mat_C_ch_6_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [0:0] m_axi_mat_C_ch_6_ARID;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [7:0] m_axi_mat_C_ch_6_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output m_axi_mat_C_ch_6_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [2:0] m_axi_mat_C_ch_6_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [3:0] m_axi_mat_C_ch_6_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.ready" *)input m_axi_mat_C_ch_6_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.data" *)output [2:0] m_axi_mat_C_ch_6_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_6_AR.valid" *)output m_axi_mat_C_ch_6_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [63:0] m_axi_mat_C_ch_6_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [1:0] m_axi_mat_C_ch_6_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [3:0] m_axi_mat_C_ch_6_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [0:0] m_axi_mat_C_ch_6_AWID;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [7:0] m_axi_mat_C_ch_6_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output m_axi_mat_C_ch_6_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [2:0] m_axi_mat_C_ch_6_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [3:0] m_axi_mat_C_ch_6_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.ready" *)input m_axi_mat_C_ch_6_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.data" *)output [2:0] m_axi_mat_C_ch_6_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_6_AW.valid" *)output m_axi_mat_C_ch_6_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_6_B.data" *)input [0:0] m_axi_mat_C_ch_6_BID;
  (* RS_HS = "m_axi_mat_C_ch_6_B.ready" *)output m_axi_mat_C_ch_6_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_6_B.data" *)input [1:0] m_axi_mat_C_ch_6_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_6_B.valid" *)input m_axi_mat_C_ch_6_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_6_R.data" *)input [511:0] m_axi_mat_C_ch_6_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_6_R.data" *)input [0:0] m_axi_mat_C_ch_6_RID;
  (* RS_HS = "m_axi_mat_C_ch_6_R.data" *)input m_axi_mat_C_ch_6_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_6_R.ready" *)output m_axi_mat_C_ch_6_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_6_R.data" *)input [1:0] m_axi_mat_C_ch_6_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_6_R.valid" *)input m_axi_mat_C_ch_6_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_6_W.data" *)output [511:0] m_axi_mat_C_ch_6_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_6_W.data" *)output m_axi_mat_C_ch_6_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_6_W.ready" *)input m_axi_mat_C_ch_6_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_6_W.data" *)output [63:0] m_axi_mat_C_ch_6_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_6_W.valid" *)output m_axi_mat_C_ch_6_WVALID;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [63:0] m_axi_mat_C_ch_7_ARADDR;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [1:0] m_axi_mat_C_ch_7_ARBURST;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [3:0] m_axi_mat_C_ch_7_ARCACHE;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [0:0] m_axi_mat_C_ch_7_ARID;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [7:0] m_axi_mat_C_ch_7_ARLEN;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output m_axi_mat_C_ch_7_ARLOCK;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [2:0] m_axi_mat_C_ch_7_ARPROT;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [3:0] m_axi_mat_C_ch_7_ARQOS;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.ready" *)input m_axi_mat_C_ch_7_ARREADY;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.data" *)output [2:0] m_axi_mat_C_ch_7_ARSIZE;
  (* RS_HS = "m_axi_mat_C_ch_7_AR.valid" *)output m_axi_mat_C_ch_7_ARVALID;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [63:0] m_axi_mat_C_ch_7_AWADDR;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [1:0] m_axi_mat_C_ch_7_AWBURST;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [3:0] m_axi_mat_C_ch_7_AWCACHE;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [0:0] m_axi_mat_C_ch_7_AWID;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [7:0] m_axi_mat_C_ch_7_AWLEN;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output m_axi_mat_C_ch_7_AWLOCK;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [2:0] m_axi_mat_C_ch_7_AWPROT;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [3:0] m_axi_mat_C_ch_7_AWQOS;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.ready" *)input m_axi_mat_C_ch_7_AWREADY;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.data" *)output [2:0] m_axi_mat_C_ch_7_AWSIZE;
  (* RS_HS = "m_axi_mat_C_ch_7_AW.valid" *)output m_axi_mat_C_ch_7_AWVALID;
  (* RS_HS = "m_axi_mat_C_ch_7_B.data" *)input [0:0] m_axi_mat_C_ch_7_BID;
  (* RS_HS = "m_axi_mat_C_ch_7_B.ready" *)output m_axi_mat_C_ch_7_BREADY;
  (* RS_HS = "m_axi_mat_C_ch_7_B.data" *)input [1:0] m_axi_mat_C_ch_7_BRESP;
  (* RS_HS = "m_axi_mat_C_ch_7_B.valid" *)input m_axi_mat_C_ch_7_BVALID;
  (* RS_HS = "m_axi_mat_C_ch_7_R.data" *)input [511:0] m_axi_mat_C_ch_7_RDATA;
  (* RS_HS = "m_axi_mat_C_ch_7_R.data" *)input [0:0] m_axi_mat_C_ch_7_RID;
  (* RS_HS = "m_axi_mat_C_ch_7_R.data" *)input m_axi_mat_C_ch_7_RLAST;
  (* RS_HS = "m_axi_mat_C_ch_7_R.ready" *)output m_axi_mat_C_ch_7_RREADY;
  (* RS_HS = "m_axi_mat_C_ch_7_R.data" *)input [1:0] m_axi_mat_C_ch_7_RRESP;
  (* RS_HS = "m_axi_mat_C_ch_7_R.valid" *)input m_axi_mat_C_ch_7_RVALID;
  (* RS_HS = "m_axi_mat_C_ch_7_W.data" *)output [511:0] m_axi_mat_C_ch_7_WDATA;
  (* RS_HS = "m_axi_mat_C_ch_7_W.data" *)output m_axi_mat_C_ch_7_WLAST;
  (* RS_HS = "m_axi_mat_C_ch_7_W.ready" *)input m_axi_mat_C_ch_7_WREADY;
  (* RS_HS = "m_axi_mat_C_ch_7_W.data" *)output [63:0] m_axi_mat_C_ch_7_WSTRB;
  (* RS_HS = "m_axi_mat_C_ch_7_W.valid" *)output m_axi_mat_C_ch_7_WVALID;
  wire ap_start;
  wire [63:0] edge_list_ptr;
  wire [63:0] edge_list_ch_0;
  wire [63:0] edge_list_ch_1;
  wire [63:0] edge_list_ch_2;
  wire [63:0] edge_list_ch_3;
  wire [63:0] edge_list_ch_4;
  wire [63:0] edge_list_ch_5;
  wire [63:0] edge_list_ch_6;
  wire [63:0] edge_list_ch_7;
  wire [63:0] mat_B_ch_0;
  wire [63:0] mat_B_ch_1;
  wire [63:0] mat_B_ch_2;
  wire [63:0] mat_B_ch_3;
  wire [63:0] mat_C_ch_in_0;
  wire [63:0] mat_C_ch_in_1;
  wire [63:0] mat_C_ch_in_2;
  wire [63:0] mat_C_ch_in_3;
  wire [63:0] mat_C_ch_in_4;
  wire [63:0] mat_C_ch_in_5;
  wire [63:0] mat_C_ch_in_6;
  wire [63:0] mat_C_ch_in_7;
  wire [63:0] mat_C_ch_0;
  wire [63:0] mat_C_ch_1;
  wire [63:0] mat_C_ch_2;
  wire [63:0] mat_C_ch_3;
  wire [63:0] mat_C_ch_4;
  wire [63:0] mat_C_ch_5;
  wire [63:0] mat_C_ch_6;
  wire [63:0] mat_C_ch_7;
  wire [31:0] NUM_ITE;
  wire [31:0] NUM_A_LEN;
  wire [31:0] M;
  wire [31:0] K;
  wire [31:0] P_N;
  wire [31:0] alpha_u;
  wire [31:0] beta_u;
  wire [32:0] PE_inst_Sextans_0__dout;
  wire PE_inst_Sextans_0__empty_n;
  wire PE_inst_Sextans_0__read;
  wire [32:0] PE_inst_Sextans_0__din;
  wire PE_inst_Sextans_0__full_n;
  wire PE_inst_Sextans_0__write;
  wire [32:0] PE_inst_Sextans_10__dout;
  wire PE_inst_Sextans_10__empty_n;
  wire PE_inst_Sextans_10__read;
  wire [32:0] PE_inst_Sextans_10__din;
  wire PE_inst_Sextans_10__full_n;
  wire PE_inst_Sextans_10__write;
  wire [32:0] PE_inst_Sextans_11__dout;
  wire PE_inst_Sextans_11__empty_n;
  wire PE_inst_Sextans_11__read;
  wire [32:0] PE_inst_Sextans_11__din;
  wire PE_inst_Sextans_11__full_n;
  wire PE_inst_Sextans_11__write;
  wire [32:0] PE_inst_Sextans_12__dout;
  wire PE_inst_Sextans_12__empty_n;
  wire PE_inst_Sextans_12__read;
  wire [32:0] PE_inst_Sextans_12__din;
  wire PE_inst_Sextans_12__full_n;
  wire PE_inst_Sextans_12__write;
  wire [32:0] PE_inst_Sextans_13__dout;
  wire PE_inst_Sextans_13__empty_n;
  wire PE_inst_Sextans_13__read;
  wire [32:0] PE_inst_Sextans_13__din;
  wire PE_inst_Sextans_13__full_n;
  wire PE_inst_Sextans_13__write;
  wire [32:0] PE_inst_Sextans_14__dout;
  wire PE_inst_Sextans_14__empty_n;
  wire PE_inst_Sextans_14__read;
  wire [32:0] PE_inst_Sextans_14__din;
  wire PE_inst_Sextans_14__full_n;
  wire PE_inst_Sextans_14__write;
  wire [32:0] PE_inst_Sextans_15__dout;
  wire PE_inst_Sextans_15__empty_n;
  wire PE_inst_Sextans_15__read;
  wire [32:0] PE_inst_Sextans_15__din;
  wire PE_inst_Sextans_15__full_n;
  wire PE_inst_Sextans_15__write;
  wire [32:0] PE_inst_Sextans_16__dout;
  wire PE_inst_Sextans_16__empty_n;
  wire PE_inst_Sextans_16__read;
  wire [32:0] PE_inst_Sextans_16__din;
  wire PE_inst_Sextans_16__full_n;
  wire PE_inst_Sextans_16__write;
  wire [32:0] PE_inst_Sextans_1__dout;
  wire PE_inst_Sextans_1__empty_n;
  wire PE_inst_Sextans_1__read;
  wire [32:0] PE_inst_Sextans_1__din;
  wire PE_inst_Sextans_1__full_n;
  wire PE_inst_Sextans_1__write;
  wire [32:0] PE_inst_Sextans_2__dout;
  wire PE_inst_Sextans_2__empty_n;
  wire PE_inst_Sextans_2__read;
  wire [32:0] PE_inst_Sextans_2__din;
  wire PE_inst_Sextans_2__full_n;
  wire PE_inst_Sextans_2__write;
  wire [32:0] PE_inst_Sextans_3__dout;
  wire PE_inst_Sextans_3__empty_n;
  wire PE_inst_Sextans_3__read;
  wire [32:0] PE_inst_Sextans_3__din;
  wire PE_inst_Sextans_3__full_n;
  wire PE_inst_Sextans_3__write;
  wire [32:0] PE_inst_Sextans_4__dout;
  wire PE_inst_Sextans_4__empty_n;
  wire PE_inst_Sextans_4__read;
  wire [32:0] PE_inst_Sextans_4__din;
  wire PE_inst_Sextans_4__full_n;
  wire PE_inst_Sextans_4__write;
  wire [32:0] PE_inst_Sextans_5__dout;
  wire PE_inst_Sextans_5__empty_n;
  wire PE_inst_Sextans_5__read;
  wire [32:0] PE_inst_Sextans_5__din;
  wire PE_inst_Sextans_5__full_n;
  wire PE_inst_Sextans_5__write;
  wire [32:0] PE_inst_Sextans_6__dout;
  wire PE_inst_Sextans_6__empty_n;
  wire PE_inst_Sextans_6__read;
  wire [32:0] PE_inst_Sextans_6__din;
  wire PE_inst_Sextans_6__full_n;
  wire PE_inst_Sextans_6__write;
  wire [32:0] PE_inst_Sextans_7__dout;
  wire PE_inst_Sextans_7__empty_n;
  wire PE_inst_Sextans_7__read;
  wire [32:0] PE_inst_Sextans_7__din;
  wire PE_inst_Sextans_7__full_n;
  wire PE_inst_Sextans_7__write;
  wire [32:0] PE_inst_Sextans_8__dout;
  wire PE_inst_Sextans_8__empty_n;
  wire PE_inst_Sextans_8__read;
  wire [32:0] PE_inst_Sextans_8__din;
  wire PE_inst_Sextans_8__full_n;
  wire PE_inst_Sextans_8__write;
  wire [32:0] PE_inst_Sextans_9__dout;
  wire PE_inst_Sextans_9__empty_n;
  wire PE_inst_Sextans_9__read;
  wire [32:0] PE_inst_Sextans_9__din;
  wire PE_inst_Sextans_9__full_n;
  wire PE_inst_Sextans_9__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_0__dout;
  wire PE_inst_to_Cmtx_Sextans_0__empty_n;
  wire PE_inst_to_Cmtx_Sextans_0__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_0__din;
  wire PE_inst_to_Cmtx_Sextans_0__full_n;
  wire PE_inst_to_Cmtx_Sextans_0__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_10__dout;
  wire PE_inst_to_Cmtx_Sextans_10__empty_n;
  wire PE_inst_to_Cmtx_Sextans_10__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_10__din;
  wire PE_inst_to_Cmtx_Sextans_10__full_n;
  wire PE_inst_to_Cmtx_Sextans_10__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_11__dout;
  wire PE_inst_to_Cmtx_Sextans_11__empty_n;
  wire PE_inst_to_Cmtx_Sextans_11__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_11__din;
  wire PE_inst_to_Cmtx_Sextans_11__full_n;
  wire PE_inst_to_Cmtx_Sextans_11__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_12__dout;
  wire PE_inst_to_Cmtx_Sextans_12__empty_n;
  wire PE_inst_to_Cmtx_Sextans_12__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_12__din;
  wire PE_inst_to_Cmtx_Sextans_12__full_n;
  wire PE_inst_to_Cmtx_Sextans_12__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_13__dout;
  wire PE_inst_to_Cmtx_Sextans_13__empty_n;
  wire PE_inst_to_Cmtx_Sextans_13__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_13__din;
  wire PE_inst_to_Cmtx_Sextans_13__full_n;
  wire PE_inst_to_Cmtx_Sextans_13__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_14__dout;
  wire PE_inst_to_Cmtx_Sextans_14__empty_n;
  wire PE_inst_to_Cmtx_Sextans_14__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_14__din;
  wire PE_inst_to_Cmtx_Sextans_14__full_n;
  wire PE_inst_to_Cmtx_Sextans_14__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_15__dout;
  wire PE_inst_to_Cmtx_Sextans_15__empty_n;
  wire PE_inst_to_Cmtx_Sextans_15__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_15__din;
  wire PE_inst_to_Cmtx_Sextans_15__full_n;
  wire PE_inst_to_Cmtx_Sextans_15__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_1__dout;
  wire PE_inst_to_Cmtx_Sextans_1__empty_n;
  wire PE_inst_to_Cmtx_Sextans_1__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_1__din;
  wire PE_inst_to_Cmtx_Sextans_1__full_n;
  wire PE_inst_to_Cmtx_Sextans_1__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_2__dout;
  wire PE_inst_to_Cmtx_Sextans_2__empty_n;
  wire PE_inst_to_Cmtx_Sextans_2__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_2__din;
  wire PE_inst_to_Cmtx_Sextans_2__full_n;
  wire PE_inst_to_Cmtx_Sextans_2__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_3__dout;
  wire PE_inst_to_Cmtx_Sextans_3__empty_n;
  wire PE_inst_to_Cmtx_Sextans_3__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_3__din;
  wire PE_inst_to_Cmtx_Sextans_3__full_n;
  wire PE_inst_to_Cmtx_Sextans_3__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_4__dout;
  wire PE_inst_to_Cmtx_Sextans_4__empty_n;
  wire PE_inst_to_Cmtx_Sextans_4__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_4__din;
  wire PE_inst_to_Cmtx_Sextans_4__full_n;
  wire PE_inst_to_Cmtx_Sextans_4__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_5__dout;
  wire PE_inst_to_Cmtx_Sextans_5__empty_n;
  wire PE_inst_to_Cmtx_Sextans_5__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_5__din;
  wire PE_inst_to_Cmtx_Sextans_5__full_n;
  wire PE_inst_to_Cmtx_Sextans_5__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_6__dout;
  wire PE_inst_to_Cmtx_Sextans_6__empty_n;
  wire PE_inst_to_Cmtx_Sextans_6__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_6__din;
  wire PE_inst_to_Cmtx_Sextans_6__full_n;
  wire PE_inst_to_Cmtx_Sextans_6__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_7__dout;
  wire PE_inst_to_Cmtx_Sextans_7__empty_n;
  wire PE_inst_to_Cmtx_Sextans_7__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_7__din;
  wire PE_inst_to_Cmtx_Sextans_7__full_n;
  wire PE_inst_to_Cmtx_Sextans_7__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_8__dout;
  wire PE_inst_to_Cmtx_Sextans_8__empty_n;
  wire PE_inst_to_Cmtx_Sextans_8__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_8__din;
  wire PE_inst_to_Cmtx_Sextans_8__full_n;
  wire PE_inst_to_Cmtx_Sextans_8__write;
  wire [32:0] PE_inst_to_Cmtx_Sextans_9__dout;
  wire PE_inst_to_Cmtx_Sextans_9__empty_n;
  wire PE_inst_to_Cmtx_Sextans_9__read;
  wire [32:0] PE_inst_to_Cmtx_Sextans_9__din;
  wire PE_inst_to_Cmtx_Sextans_9__full_n;
  wire PE_inst_to_Cmtx_Sextans_9__write;
  wire [512:0] fifo_A_Sextans_0__dout;
  wire fifo_A_Sextans_0__empty_n;
  wire fifo_A_Sextans_0__read;
  wire [512:0] fifo_A_Sextans_0__din;
  wire fifo_A_Sextans_0__full_n;
  wire fifo_A_Sextans_0__write;
  wire [512:0] fifo_A_Sextans_1__dout;
  wire fifo_A_Sextans_1__empty_n;
  wire fifo_A_Sextans_1__read;
  wire [512:0] fifo_A_Sextans_1__din;
  wire fifo_A_Sextans_1__full_n;
  wire fifo_A_Sextans_1__write;
  wire [512:0] fifo_A_Sextans_2__dout;
  wire fifo_A_Sextans_2__empty_n;
  wire fifo_A_Sextans_2__read;
  wire [512:0] fifo_A_Sextans_2__din;
  wire fifo_A_Sextans_2__full_n;
  wire fifo_A_Sextans_2__write;
  wire [512:0] fifo_A_Sextans_3__dout;
  wire fifo_A_Sextans_3__empty_n;
  wire fifo_A_Sextans_3__read;
  wire [512:0] fifo_A_Sextans_3__din;
  wire fifo_A_Sextans_3__full_n;
  wire fifo_A_Sextans_3__write;
  wire [512:0] fifo_A_Sextans_4__dout;
  wire fifo_A_Sextans_4__empty_n;
  wire fifo_A_Sextans_4__read;
  wire [512:0] fifo_A_Sextans_4__din;
  wire fifo_A_Sextans_4__full_n;
  wire fifo_A_Sextans_4__write;
  wire [512:0] fifo_A_Sextans_5__dout;
  wire fifo_A_Sextans_5__empty_n;
  wire fifo_A_Sextans_5__read;
  wire [512:0] fifo_A_Sextans_5__din;
  wire fifo_A_Sextans_5__full_n;
  wire fifo_A_Sextans_5__write;
  wire [512:0] fifo_A_Sextans_6__dout;
  wire fifo_A_Sextans_6__empty_n;
  wire fifo_A_Sextans_6__read;
  wire [512:0] fifo_A_Sextans_6__din;
  wire fifo_A_Sextans_6__full_n;
  wire fifo_A_Sextans_6__write;
  wire [512:0] fifo_A_Sextans_7__dout;
  wire fifo_A_Sextans_7__empty_n;
  wire fifo_A_Sextans_7__read;
  wire [512:0] fifo_A_Sextans_7__din;
  wire fifo_A_Sextans_7__full_n;
  wire fifo_A_Sextans_7__write;
  wire [256:0] fifo_A_pe_Sextans_0__dout;
  wire fifo_A_pe_Sextans_0__empty_n;
  wire fifo_A_pe_Sextans_0__read;
  wire [256:0] fifo_A_pe_Sextans_0__din;
  wire fifo_A_pe_Sextans_0__full_n;
  wire fifo_A_pe_Sextans_0__write;
  wire [256:0] fifo_A_pe_Sextans_10__dout;
  wire fifo_A_pe_Sextans_10__empty_n;
  wire fifo_A_pe_Sextans_10__read;
  wire [256:0] fifo_A_pe_Sextans_10__din;
  wire fifo_A_pe_Sextans_10__full_n;
  wire fifo_A_pe_Sextans_10__write;
  wire [256:0] fifo_A_pe_Sextans_11__dout;
  wire fifo_A_pe_Sextans_11__empty_n;
  wire fifo_A_pe_Sextans_11__read;
  wire [256:0] fifo_A_pe_Sextans_11__din;
  wire fifo_A_pe_Sextans_11__full_n;
  wire fifo_A_pe_Sextans_11__write;
  wire [256:0] fifo_A_pe_Sextans_12__dout;
  wire fifo_A_pe_Sextans_12__empty_n;
  wire fifo_A_pe_Sextans_12__read;
  wire [256:0] fifo_A_pe_Sextans_12__din;
  wire fifo_A_pe_Sextans_12__full_n;
  wire fifo_A_pe_Sextans_12__write;
  wire [256:0] fifo_A_pe_Sextans_13__dout;
  wire fifo_A_pe_Sextans_13__empty_n;
  wire fifo_A_pe_Sextans_13__read;
  wire [256:0] fifo_A_pe_Sextans_13__din;
  wire fifo_A_pe_Sextans_13__full_n;
  wire fifo_A_pe_Sextans_13__write;
  wire [256:0] fifo_A_pe_Sextans_14__dout;
  wire fifo_A_pe_Sextans_14__empty_n;
  wire fifo_A_pe_Sextans_14__read;
  wire [256:0] fifo_A_pe_Sextans_14__din;
  wire fifo_A_pe_Sextans_14__full_n;
  wire fifo_A_pe_Sextans_14__write;
  wire [256:0] fifo_A_pe_Sextans_15__dout;
  wire fifo_A_pe_Sextans_15__empty_n;
  wire fifo_A_pe_Sextans_15__read;
  wire [256:0] fifo_A_pe_Sextans_15__din;
  wire fifo_A_pe_Sextans_15__full_n;
  wire fifo_A_pe_Sextans_15__write;
  wire [256:0] fifo_A_pe_Sextans_1__dout;
  wire fifo_A_pe_Sextans_1__empty_n;
  wire fifo_A_pe_Sextans_1__read;
  wire [256:0] fifo_A_pe_Sextans_1__din;
  wire fifo_A_pe_Sextans_1__full_n;
  wire fifo_A_pe_Sextans_1__write;
  wire [256:0] fifo_A_pe_Sextans_2__dout;
  wire fifo_A_pe_Sextans_2__empty_n;
  wire fifo_A_pe_Sextans_2__read;
  wire [256:0] fifo_A_pe_Sextans_2__din;
  wire fifo_A_pe_Sextans_2__full_n;
  wire fifo_A_pe_Sextans_2__write;
  wire [256:0] fifo_A_pe_Sextans_3__dout;
  wire fifo_A_pe_Sextans_3__empty_n;
  wire fifo_A_pe_Sextans_3__read;
  wire [256:0] fifo_A_pe_Sextans_3__din;
  wire fifo_A_pe_Sextans_3__full_n;
  wire fifo_A_pe_Sextans_3__write;
  wire [256:0] fifo_A_pe_Sextans_4__dout;
  wire fifo_A_pe_Sextans_4__empty_n;
  wire fifo_A_pe_Sextans_4__read;
  wire [256:0] fifo_A_pe_Sextans_4__din;
  wire fifo_A_pe_Sextans_4__full_n;
  wire fifo_A_pe_Sextans_4__write;
  wire [256:0] fifo_A_pe_Sextans_5__dout;
  wire fifo_A_pe_Sextans_5__empty_n;
  wire fifo_A_pe_Sextans_5__read;
  wire [256:0] fifo_A_pe_Sextans_5__din;
  wire fifo_A_pe_Sextans_5__full_n;
  wire fifo_A_pe_Sextans_5__write;
  wire [256:0] fifo_A_pe_Sextans_6__dout;
  wire fifo_A_pe_Sextans_6__empty_n;
  wire fifo_A_pe_Sextans_6__read;
  wire [256:0] fifo_A_pe_Sextans_6__din;
  wire fifo_A_pe_Sextans_6__full_n;
  wire fifo_A_pe_Sextans_6__write;
  wire [256:0] fifo_A_pe_Sextans_7__dout;
  wire fifo_A_pe_Sextans_7__empty_n;
  wire fifo_A_pe_Sextans_7__read;
  wire [256:0] fifo_A_pe_Sextans_7__din;
  wire fifo_A_pe_Sextans_7__full_n;
  wire fifo_A_pe_Sextans_7__write;
  wire [256:0] fifo_A_pe_Sextans_8__dout;
  wire fifo_A_pe_Sextans_8__empty_n;
  wire fifo_A_pe_Sextans_8__read;
  wire [256:0] fifo_A_pe_Sextans_8__din;
  wire fifo_A_pe_Sextans_8__full_n;
  wire fifo_A_pe_Sextans_8__write;
  wire [256:0] fifo_A_pe_Sextans_9__dout;
  wire fifo_A_pe_Sextans_9__empty_n;
  wire fifo_A_pe_Sextans_9__read;
  wire [256:0] fifo_A_pe_Sextans_9__din;
  wire fifo_A_pe_Sextans_9__full_n;
  wire fifo_A_pe_Sextans_9__write;
  wire [512:0] fifo_B_pe_Sextans_0__dout;
  wire fifo_B_pe_Sextans_0__empty_n;
  wire fifo_B_pe_Sextans_0__read;
  wire [512:0] fifo_B_pe_Sextans_0__din;
  wire fifo_B_pe_Sextans_0__full_n;
  wire fifo_B_pe_Sextans_0__write;
  wire [512:0] fifo_B_pe_Sextans_10__dout;
  wire fifo_B_pe_Sextans_10__empty_n;
  wire fifo_B_pe_Sextans_10__read;
  wire [512:0] fifo_B_pe_Sextans_10__din;
  wire fifo_B_pe_Sextans_10__full_n;
  wire fifo_B_pe_Sextans_10__write;
  wire [512:0] fifo_B_pe_Sextans_11__dout;
  wire fifo_B_pe_Sextans_11__empty_n;
  wire fifo_B_pe_Sextans_11__read;
  wire [512:0] fifo_B_pe_Sextans_11__din;
  wire fifo_B_pe_Sextans_11__full_n;
  wire fifo_B_pe_Sextans_11__write;
  wire [512:0] fifo_B_pe_Sextans_12__dout;
  wire fifo_B_pe_Sextans_12__empty_n;
  wire fifo_B_pe_Sextans_12__read;
  wire [512:0] fifo_B_pe_Sextans_12__din;
  wire fifo_B_pe_Sextans_12__full_n;
  wire fifo_B_pe_Sextans_12__write;
  wire [512:0] fifo_B_pe_Sextans_13__dout;
  wire fifo_B_pe_Sextans_13__empty_n;
  wire fifo_B_pe_Sextans_13__read;
  wire [512:0] fifo_B_pe_Sextans_13__din;
  wire fifo_B_pe_Sextans_13__full_n;
  wire fifo_B_pe_Sextans_13__write;
  wire [512:0] fifo_B_pe_Sextans_14__dout;
  wire fifo_B_pe_Sextans_14__empty_n;
  wire fifo_B_pe_Sextans_14__read;
  wire [512:0] fifo_B_pe_Sextans_14__din;
  wire fifo_B_pe_Sextans_14__full_n;
  wire fifo_B_pe_Sextans_14__write;
  wire [512:0] fifo_B_pe_Sextans_15__dout;
  wire fifo_B_pe_Sextans_15__empty_n;
  wire fifo_B_pe_Sextans_15__read;
  wire [512:0] fifo_B_pe_Sextans_15__din;
  wire fifo_B_pe_Sextans_15__full_n;
  wire fifo_B_pe_Sextans_15__write;
  wire [512:0] fifo_B_pe_Sextans_16__dout;
  wire fifo_B_pe_Sextans_16__empty_n;
  wire fifo_B_pe_Sextans_16__read;
  wire [512:0] fifo_B_pe_Sextans_16__din;
  wire fifo_B_pe_Sextans_16__full_n;
  wire fifo_B_pe_Sextans_16__write;
  wire [512:0] fifo_B_pe_Sextans_17__dout;
  wire fifo_B_pe_Sextans_17__empty_n;
  wire fifo_B_pe_Sextans_17__read;
  wire [512:0] fifo_B_pe_Sextans_17__din;
  wire fifo_B_pe_Sextans_17__full_n;
  wire fifo_B_pe_Sextans_17__write;
  wire [512:0] fifo_B_pe_Sextans_18__dout;
  wire fifo_B_pe_Sextans_18__empty_n;
  wire fifo_B_pe_Sextans_18__read;
  wire [512:0] fifo_B_pe_Sextans_18__din;
  wire fifo_B_pe_Sextans_18__full_n;
  wire fifo_B_pe_Sextans_18__write;
  wire [512:0] fifo_B_pe_Sextans_19__dout;
  wire fifo_B_pe_Sextans_19__empty_n;
  wire fifo_B_pe_Sextans_19__read;
  wire [512:0] fifo_B_pe_Sextans_19__din;
  wire fifo_B_pe_Sextans_19__full_n;
  wire fifo_B_pe_Sextans_19__write;
  wire [512:0] fifo_B_pe_Sextans_1__dout;
  wire fifo_B_pe_Sextans_1__empty_n;
  wire fifo_B_pe_Sextans_1__read;
  wire [512:0] fifo_B_pe_Sextans_1__din;
  wire fifo_B_pe_Sextans_1__full_n;
  wire fifo_B_pe_Sextans_1__write;
  wire [512:0] fifo_B_pe_Sextans_20__dout;
  wire fifo_B_pe_Sextans_20__empty_n;
  wire fifo_B_pe_Sextans_20__read;
  wire [512:0] fifo_B_pe_Sextans_20__din;
  wire fifo_B_pe_Sextans_20__full_n;
  wire fifo_B_pe_Sextans_20__write;
  wire [512:0] fifo_B_pe_Sextans_21__dout;
  wire fifo_B_pe_Sextans_21__empty_n;
  wire fifo_B_pe_Sextans_21__read;
  wire [512:0] fifo_B_pe_Sextans_21__din;
  wire fifo_B_pe_Sextans_21__full_n;
  wire fifo_B_pe_Sextans_21__write;
  wire [512:0] fifo_B_pe_Sextans_22__dout;
  wire fifo_B_pe_Sextans_22__empty_n;
  wire fifo_B_pe_Sextans_22__read;
  wire [512:0] fifo_B_pe_Sextans_22__din;
  wire fifo_B_pe_Sextans_22__full_n;
  wire fifo_B_pe_Sextans_22__write;
  wire [512:0] fifo_B_pe_Sextans_23__dout;
  wire fifo_B_pe_Sextans_23__empty_n;
  wire fifo_B_pe_Sextans_23__read;
  wire [512:0] fifo_B_pe_Sextans_23__din;
  wire fifo_B_pe_Sextans_23__full_n;
  wire fifo_B_pe_Sextans_23__write;
  wire [512:0] fifo_B_pe_Sextans_24__dout;
  wire fifo_B_pe_Sextans_24__empty_n;
  wire fifo_B_pe_Sextans_24__read;
  wire [512:0] fifo_B_pe_Sextans_24__din;
  wire fifo_B_pe_Sextans_24__full_n;
  wire fifo_B_pe_Sextans_24__write;
  wire [512:0] fifo_B_pe_Sextans_25__dout;
  wire fifo_B_pe_Sextans_25__empty_n;
  wire fifo_B_pe_Sextans_25__read;
  wire [512:0] fifo_B_pe_Sextans_25__din;
  wire fifo_B_pe_Sextans_25__full_n;
  wire fifo_B_pe_Sextans_25__write;
  wire [512:0] fifo_B_pe_Sextans_26__dout;
  wire fifo_B_pe_Sextans_26__empty_n;
  wire fifo_B_pe_Sextans_26__read;
  wire [512:0] fifo_B_pe_Sextans_26__din;
  wire fifo_B_pe_Sextans_26__full_n;
  wire fifo_B_pe_Sextans_26__write;
  wire [512:0] fifo_B_pe_Sextans_27__dout;
  wire fifo_B_pe_Sextans_27__empty_n;
  wire fifo_B_pe_Sextans_27__read;
  wire [512:0] fifo_B_pe_Sextans_27__din;
  wire fifo_B_pe_Sextans_27__full_n;
  wire fifo_B_pe_Sextans_27__write;
  wire [512:0] fifo_B_pe_Sextans_28__dout;
  wire fifo_B_pe_Sextans_28__empty_n;
  wire fifo_B_pe_Sextans_28__read;
  wire [512:0] fifo_B_pe_Sextans_28__din;
  wire fifo_B_pe_Sextans_28__full_n;
  wire fifo_B_pe_Sextans_28__write;
  wire [512:0] fifo_B_pe_Sextans_29__dout;
  wire fifo_B_pe_Sextans_29__empty_n;
  wire fifo_B_pe_Sextans_29__read;
  wire [512:0] fifo_B_pe_Sextans_29__din;
  wire fifo_B_pe_Sextans_29__full_n;
  wire fifo_B_pe_Sextans_29__write;
  wire [512:0] fifo_B_pe_Sextans_2__dout;
  wire fifo_B_pe_Sextans_2__empty_n;
  wire fifo_B_pe_Sextans_2__read;
  wire [512:0] fifo_B_pe_Sextans_2__din;
  wire fifo_B_pe_Sextans_2__full_n;
  wire fifo_B_pe_Sextans_2__write;
  wire [512:0] fifo_B_pe_Sextans_30__dout;
  wire fifo_B_pe_Sextans_30__empty_n;
  wire fifo_B_pe_Sextans_30__read;
  wire [512:0] fifo_B_pe_Sextans_30__din;
  wire fifo_B_pe_Sextans_30__full_n;
  wire fifo_B_pe_Sextans_30__write;
  wire [512:0] fifo_B_pe_Sextans_31__dout;
  wire fifo_B_pe_Sextans_31__empty_n;
  wire fifo_B_pe_Sextans_31__read;
  wire [512:0] fifo_B_pe_Sextans_31__din;
  wire fifo_B_pe_Sextans_31__full_n;
  wire fifo_B_pe_Sextans_31__write;
  wire [512:0] fifo_B_pe_Sextans_32__dout;
  wire fifo_B_pe_Sextans_32__empty_n;
  wire fifo_B_pe_Sextans_32__read;
  wire [512:0] fifo_B_pe_Sextans_32__din;
  wire fifo_B_pe_Sextans_32__full_n;
  wire fifo_B_pe_Sextans_32__write;
  wire [512:0] fifo_B_pe_Sextans_33__dout;
  wire fifo_B_pe_Sextans_33__empty_n;
  wire fifo_B_pe_Sextans_33__read;
  wire [512:0] fifo_B_pe_Sextans_33__din;
  wire fifo_B_pe_Sextans_33__full_n;
  wire fifo_B_pe_Sextans_33__write;
  wire [512:0] fifo_B_pe_Sextans_34__dout;
  wire fifo_B_pe_Sextans_34__empty_n;
  wire fifo_B_pe_Sextans_34__read;
  wire [512:0] fifo_B_pe_Sextans_34__din;
  wire fifo_B_pe_Sextans_34__full_n;
  wire fifo_B_pe_Sextans_34__write;
  wire [512:0] fifo_B_pe_Sextans_35__dout;
  wire fifo_B_pe_Sextans_35__empty_n;
  wire fifo_B_pe_Sextans_35__read;
  wire [512:0] fifo_B_pe_Sextans_35__din;
  wire fifo_B_pe_Sextans_35__full_n;
  wire fifo_B_pe_Sextans_35__write;
  wire [512:0] fifo_B_pe_Sextans_36__dout;
  wire fifo_B_pe_Sextans_36__empty_n;
  wire fifo_B_pe_Sextans_36__read;
  wire [512:0] fifo_B_pe_Sextans_36__din;
  wire fifo_B_pe_Sextans_36__full_n;
  wire fifo_B_pe_Sextans_36__write;
  wire [512:0] fifo_B_pe_Sextans_37__dout;
  wire fifo_B_pe_Sextans_37__empty_n;
  wire fifo_B_pe_Sextans_37__read;
  wire [512:0] fifo_B_pe_Sextans_37__din;
  wire fifo_B_pe_Sextans_37__full_n;
  wire fifo_B_pe_Sextans_37__write;
  wire [512:0] fifo_B_pe_Sextans_38__dout;
  wire fifo_B_pe_Sextans_38__empty_n;
  wire fifo_B_pe_Sextans_38__read;
  wire [512:0] fifo_B_pe_Sextans_38__din;
  wire fifo_B_pe_Sextans_38__full_n;
  wire fifo_B_pe_Sextans_38__write;
  wire [512:0] fifo_B_pe_Sextans_39__dout;
  wire fifo_B_pe_Sextans_39__empty_n;
  wire fifo_B_pe_Sextans_39__read;
  wire [512:0] fifo_B_pe_Sextans_39__din;
  wire fifo_B_pe_Sextans_39__full_n;
  wire fifo_B_pe_Sextans_39__write;
  wire [512:0] fifo_B_pe_Sextans_3__dout;
  wire fifo_B_pe_Sextans_3__empty_n;
  wire fifo_B_pe_Sextans_3__read;
  wire [512:0] fifo_B_pe_Sextans_3__din;
  wire fifo_B_pe_Sextans_3__full_n;
  wire fifo_B_pe_Sextans_3__write;
  wire [512:0] fifo_B_pe_Sextans_40__dout;
  wire fifo_B_pe_Sextans_40__empty_n;
  wire fifo_B_pe_Sextans_40__read;
  wire [512:0] fifo_B_pe_Sextans_40__din;
  wire fifo_B_pe_Sextans_40__full_n;
  wire fifo_B_pe_Sextans_40__write;
  wire [512:0] fifo_B_pe_Sextans_41__dout;
  wire fifo_B_pe_Sextans_41__empty_n;
  wire fifo_B_pe_Sextans_41__read;
  wire [512:0] fifo_B_pe_Sextans_41__din;
  wire fifo_B_pe_Sextans_41__full_n;
  wire fifo_B_pe_Sextans_41__write;
  wire [512:0] fifo_B_pe_Sextans_42__dout;
  wire fifo_B_pe_Sextans_42__empty_n;
  wire fifo_B_pe_Sextans_42__read;
  wire [512:0] fifo_B_pe_Sextans_42__din;
  wire fifo_B_pe_Sextans_42__full_n;
  wire fifo_B_pe_Sextans_42__write;
  wire [512:0] fifo_B_pe_Sextans_43__dout;
  wire fifo_B_pe_Sextans_43__empty_n;
  wire fifo_B_pe_Sextans_43__read;
  wire [512:0] fifo_B_pe_Sextans_43__din;
  wire fifo_B_pe_Sextans_43__full_n;
  wire fifo_B_pe_Sextans_43__write;
  wire [512:0] fifo_B_pe_Sextans_44__dout;
  wire fifo_B_pe_Sextans_44__empty_n;
  wire fifo_B_pe_Sextans_44__read;
  wire [512:0] fifo_B_pe_Sextans_44__din;
  wire fifo_B_pe_Sextans_44__full_n;
  wire fifo_B_pe_Sextans_44__write;
  wire [512:0] fifo_B_pe_Sextans_45__dout;
  wire fifo_B_pe_Sextans_45__empty_n;
  wire fifo_B_pe_Sextans_45__read;
  wire [512:0] fifo_B_pe_Sextans_45__din;
  wire fifo_B_pe_Sextans_45__full_n;
  wire fifo_B_pe_Sextans_45__write;
  wire [512:0] fifo_B_pe_Sextans_46__dout;
  wire fifo_B_pe_Sextans_46__empty_n;
  wire fifo_B_pe_Sextans_46__read;
  wire [512:0] fifo_B_pe_Sextans_46__din;
  wire fifo_B_pe_Sextans_46__full_n;
  wire fifo_B_pe_Sextans_46__write;
  wire [512:0] fifo_B_pe_Sextans_47__dout;
  wire fifo_B_pe_Sextans_47__empty_n;
  wire fifo_B_pe_Sextans_47__read;
  wire [512:0] fifo_B_pe_Sextans_47__din;
  wire fifo_B_pe_Sextans_47__full_n;
  wire fifo_B_pe_Sextans_47__write;
  wire [512:0] fifo_B_pe_Sextans_48__dout;
  wire fifo_B_pe_Sextans_48__empty_n;
  wire fifo_B_pe_Sextans_48__read;
  wire [512:0] fifo_B_pe_Sextans_48__din;
  wire fifo_B_pe_Sextans_48__full_n;
  wire fifo_B_pe_Sextans_48__write;
  wire [512:0] fifo_B_pe_Sextans_49__dout;
  wire fifo_B_pe_Sextans_49__empty_n;
  wire fifo_B_pe_Sextans_49__read;
  wire [512:0] fifo_B_pe_Sextans_49__din;
  wire fifo_B_pe_Sextans_49__full_n;
  wire fifo_B_pe_Sextans_49__write;
  wire [512:0] fifo_B_pe_Sextans_4__dout;
  wire fifo_B_pe_Sextans_4__empty_n;
  wire fifo_B_pe_Sextans_4__read;
  wire [512:0] fifo_B_pe_Sextans_4__din;
  wire fifo_B_pe_Sextans_4__full_n;
  wire fifo_B_pe_Sextans_4__write;
  wire [512:0] fifo_B_pe_Sextans_50__dout;
  wire fifo_B_pe_Sextans_50__empty_n;
  wire fifo_B_pe_Sextans_50__read;
  wire [512:0] fifo_B_pe_Sextans_50__din;
  wire fifo_B_pe_Sextans_50__full_n;
  wire fifo_B_pe_Sextans_50__write;
  wire [512:0] fifo_B_pe_Sextans_51__dout;
  wire fifo_B_pe_Sextans_51__empty_n;
  wire fifo_B_pe_Sextans_51__read;
  wire [512:0] fifo_B_pe_Sextans_51__din;
  wire fifo_B_pe_Sextans_51__full_n;
  wire fifo_B_pe_Sextans_51__write;
  wire [512:0] fifo_B_pe_Sextans_52__dout;
  wire fifo_B_pe_Sextans_52__empty_n;
  wire fifo_B_pe_Sextans_52__read;
  wire [512:0] fifo_B_pe_Sextans_52__din;
  wire fifo_B_pe_Sextans_52__full_n;
  wire fifo_B_pe_Sextans_52__write;
  wire [512:0] fifo_B_pe_Sextans_53__dout;
  wire fifo_B_pe_Sextans_53__empty_n;
  wire fifo_B_pe_Sextans_53__read;
  wire [512:0] fifo_B_pe_Sextans_53__din;
  wire fifo_B_pe_Sextans_53__full_n;
  wire fifo_B_pe_Sextans_53__write;
  wire [512:0] fifo_B_pe_Sextans_54__dout;
  wire fifo_B_pe_Sextans_54__empty_n;
  wire fifo_B_pe_Sextans_54__read;
  wire [512:0] fifo_B_pe_Sextans_54__din;
  wire fifo_B_pe_Sextans_54__full_n;
  wire fifo_B_pe_Sextans_54__write;
  wire [512:0] fifo_B_pe_Sextans_55__dout;
  wire fifo_B_pe_Sextans_55__empty_n;
  wire fifo_B_pe_Sextans_55__read;
  wire [512:0] fifo_B_pe_Sextans_55__din;
  wire fifo_B_pe_Sextans_55__full_n;
  wire fifo_B_pe_Sextans_55__write;
  wire [512:0] fifo_B_pe_Sextans_56__dout;
  wire fifo_B_pe_Sextans_56__empty_n;
  wire fifo_B_pe_Sextans_56__read;
  wire [512:0] fifo_B_pe_Sextans_56__din;
  wire fifo_B_pe_Sextans_56__full_n;
  wire fifo_B_pe_Sextans_56__write;
  wire [512:0] fifo_B_pe_Sextans_57__dout;
  wire fifo_B_pe_Sextans_57__empty_n;
  wire fifo_B_pe_Sextans_57__read;
  wire [512:0] fifo_B_pe_Sextans_57__din;
  wire fifo_B_pe_Sextans_57__full_n;
  wire fifo_B_pe_Sextans_57__write;
  wire [512:0] fifo_B_pe_Sextans_58__dout;
  wire fifo_B_pe_Sextans_58__empty_n;
  wire fifo_B_pe_Sextans_58__read;
  wire [512:0] fifo_B_pe_Sextans_58__din;
  wire fifo_B_pe_Sextans_58__full_n;
  wire fifo_B_pe_Sextans_58__write;
  wire [512:0] fifo_B_pe_Sextans_59__dout;
  wire fifo_B_pe_Sextans_59__empty_n;
  wire fifo_B_pe_Sextans_59__read;
  wire [512:0] fifo_B_pe_Sextans_59__din;
  wire fifo_B_pe_Sextans_59__full_n;
  wire fifo_B_pe_Sextans_59__write;
  wire [512:0] fifo_B_pe_Sextans_5__dout;
  wire fifo_B_pe_Sextans_5__empty_n;
  wire fifo_B_pe_Sextans_5__read;
  wire [512:0] fifo_B_pe_Sextans_5__din;
  wire fifo_B_pe_Sextans_5__full_n;
  wire fifo_B_pe_Sextans_5__write;
  wire [512:0] fifo_B_pe_Sextans_60__dout;
  wire fifo_B_pe_Sextans_60__empty_n;
  wire fifo_B_pe_Sextans_60__read;
  wire [512:0] fifo_B_pe_Sextans_60__din;
  wire fifo_B_pe_Sextans_60__full_n;
  wire fifo_B_pe_Sextans_60__write;
  wire [512:0] fifo_B_pe_Sextans_61__dout;
  wire fifo_B_pe_Sextans_61__empty_n;
  wire fifo_B_pe_Sextans_61__read;
  wire [512:0] fifo_B_pe_Sextans_61__din;
  wire fifo_B_pe_Sextans_61__full_n;
  wire fifo_B_pe_Sextans_61__write;
  wire [512:0] fifo_B_pe_Sextans_62__dout;
  wire fifo_B_pe_Sextans_62__empty_n;
  wire fifo_B_pe_Sextans_62__read;
  wire [512:0] fifo_B_pe_Sextans_62__din;
  wire fifo_B_pe_Sextans_62__full_n;
  wire fifo_B_pe_Sextans_62__write;
  wire [512:0] fifo_B_pe_Sextans_63__dout;
  wire fifo_B_pe_Sextans_63__empty_n;
  wire fifo_B_pe_Sextans_63__read;
  wire [512:0] fifo_B_pe_Sextans_63__din;
  wire fifo_B_pe_Sextans_63__full_n;
  wire fifo_B_pe_Sextans_63__write;
  wire [512:0] fifo_B_pe_Sextans_64__dout;
  wire fifo_B_pe_Sextans_64__empty_n;
  wire fifo_B_pe_Sextans_64__read;
  wire [512:0] fifo_B_pe_Sextans_64__din;
  wire fifo_B_pe_Sextans_64__full_n;
  wire fifo_B_pe_Sextans_64__write;
  wire [512:0] fifo_B_pe_Sextans_65__dout;
  wire fifo_B_pe_Sextans_65__empty_n;
  wire fifo_B_pe_Sextans_65__read;
  wire [512:0] fifo_B_pe_Sextans_65__din;
  wire fifo_B_pe_Sextans_65__full_n;
  wire fifo_B_pe_Sextans_65__write;
  wire [512:0] fifo_B_pe_Sextans_66__dout;
  wire fifo_B_pe_Sextans_66__empty_n;
  wire fifo_B_pe_Sextans_66__read;
  wire [512:0] fifo_B_pe_Sextans_66__din;
  wire fifo_B_pe_Sextans_66__full_n;
  wire fifo_B_pe_Sextans_66__write;
  wire [512:0] fifo_B_pe_Sextans_67__dout;
  wire fifo_B_pe_Sextans_67__empty_n;
  wire fifo_B_pe_Sextans_67__read;
  wire [512:0] fifo_B_pe_Sextans_67__din;
  wire fifo_B_pe_Sextans_67__full_n;
  wire fifo_B_pe_Sextans_67__write;
  wire [512:0] fifo_B_pe_Sextans_6__dout;
  wire fifo_B_pe_Sextans_6__empty_n;
  wire fifo_B_pe_Sextans_6__read;
  wire [512:0] fifo_B_pe_Sextans_6__din;
  wire fifo_B_pe_Sextans_6__full_n;
  wire fifo_B_pe_Sextans_6__write;
  wire [512:0] fifo_B_pe_Sextans_7__dout;
  wire fifo_B_pe_Sextans_7__empty_n;
  wire fifo_B_pe_Sextans_7__read;
  wire [512:0] fifo_B_pe_Sextans_7__din;
  wire fifo_B_pe_Sextans_7__full_n;
  wire fifo_B_pe_Sextans_7__write;
  wire [512:0] fifo_B_pe_Sextans_8__dout;
  wire fifo_B_pe_Sextans_8__empty_n;
  wire fifo_B_pe_Sextans_8__read;
  wire [512:0] fifo_B_pe_Sextans_8__din;
  wire fifo_B_pe_Sextans_8__full_n;
  wire fifo_B_pe_Sextans_8__write;
  wire [512:0] fifo_B_pe_Sextans_9__dout;
  wire fifo_B_pe_Sextans_9__empty_n;
  wire fifo_B_pe_Sextans_9__read;
  wire [512:0] fifo_B_pe_Sextans_9__din;
  wire fifo_B_pe_Sextans_9__full_n;
  wire fifo_B_pe_Sextans_9__write;
  wire [512:0] fifo_C_ch_Sextans_0__dout;
  wire fifo_C_ch_Sextans_0__empty_n;
  wire fifo_C_ch_Sextans_0__read;
  wire [512:0] fifo_C_ch_Sextans_0__din;
  wire fifo_C_ch_Sextans_0__full_n;
  wire fifo_C_ch_Sextans_0__write;
  wire [512:0] fifo_C_ch_Sextans_1__dout;
  wire fifo_C_ch_Sextans_1__empty_n;
  wire fifo_C_ch_Sextans_1__read;
  wire [512:0] fifo_C_ch_Sextans_1__din;
  wire fifo_C_ch_Sextans_1__full_n;
  wire fifo_C_ch_Sextans_1__write;
  wire [512:0] fifo_C_ch_Sextans_2__dout;
  wire fifo_C_ch_Sextans_2__empty_n;
  wire fifo_C_ch_Sextans_2__read;
  wire [512:0] fifo_C_ch_Sextans_2__din;
  wire fifo_C_ch_Sextans_2__full_n;
  wire fifo_C_ch_Sextans_2__write;
  wire [512:0] fifo_C_ch_Sextans_3__dout;
  wire fifo_C_ch_Sextans_3__empty_n;
  wire fifo_C_ch_Sextans_3__read;
  wire [512:0] fifo_C_ch_Sextans_3__din;
  wire fifo_C_ch_Sextans_3__full_n;
  wire fifo_C_ch_Sextans_3__write;
  wire [512:0] fifo_C_ch_Sextans_4__dout;
  wire fifo_C_ch_Sextans_4__empty_n;
  wire fifo_C_ch_Sextans_4__read;
  wire [512:0] fifo_C_ch_Sextans_4__din;
  wire fifo_C_ch_Sextans_4__full_n;
  wire fifo_C_ch_Sextans_4__write;
  wire [512:0] fifo_C_ch_Sextans_5__dout;
  wire fifo_C_ch_Sextans_5__empty_n;
  wire fifo_C_ch_Sextans_5__read;
  wire [512:0] fifo_C_ch_Sextans_5__din;
  wire fifo_C_ch_Sextans_5__full_n;
  wire fifo_C_ch_Sextans_5__write;
  wire [512:0] fifo_C_ch_Sextans_6__dout;
  wire fifo_C_ch_Sextans_6__empty_n;
  wire fifo_C_ch_Sextans_6__read;
  wire [512:0] fifo_C_ch_Sextans_6__din;
  wire fifo_C_ch_Sextans_6__full_n;
  wire fifo_C_ch_Sextans_6__write;
  wire [512:0] fifo_C_ch_Sextans_7__dout;
  wire fifo_C_ch_Sextans_7__empty_n;
  wire fifo_C_ch_Sextans_7__read;
  wire [512:0] fifo_C_ch_Sextans_7__din;
  wire fifo_C_ch_Sextans_7__full_n;
  wire fifo_C_ch_Sextans_7__write;
  wire [512:0] fifo_C_ch_result_Sextans_0__dout;
  wire fifo_C_ch_result_Sextans_0__empty_n;
  wire fifo_C_ch_result_Sextans_0__read;
  wire [512:0] fifo_C_ch_result_Sextans_0__din;
  wire fifo_C_ch_result_Sextans_0__full_n;
  wire fifo_C_ch_result_Sextans_0__write;
  wire [512:0] fifo_C_ch_result_Sextans_1__dout;
  wire fifo_C_ch_result_Sextans_1__empty_n;
  wire fifo_C_ch_result_Sextans_1__read;
  wire [512:0] fifo_C_ch_result_Sextans_1__din;
  wire fifo_C_ch_result_Sextans_1__full_n;
  wire fifo_C_ch_result_Sextans_1__write;
  wire [512:0] fifo_C_ch_result_Sextans_2__dout;
  wire fifo_C_ch_result_Sextans_2__empty_n;
  wire fifo_C_ch_result_Sextans_2__read;
  wire [512:0] fifo_C_ch_result_Sextans_2__din;
  wire fifo_C_ch_result_Sextans_2__full_n;
  wire fifo_C_ch_result_Sextans_2__write;
  wire [512:0] fifo_C_ch_result_Sextans_3__dout;
  wire fifo_C_ch_result_Sextans_3__empty_n;
  wire fifo_C_ch_result_Sextans_3__read;
  wire [512:0] fifo_C_ch_result_Sextans_3__din;
  wire fifo_C_ch_result_Sextans_3__full_n;
  wire fifo_C_ch_result_Sextans_3__write;
  wire [512:0] fifo_C_ch_result_Sextans_4__dout;
  wire fifo_C_ch_result_Sextans_4__empty_n;
  wire fifo_C_ch_result_Sextans_4__read;
  wire [512:0] fifo_C_ch_result_Sextans_4__din;
  wire fifo_C_ch_result_Sextans_4__full_n;
  wire fifo_C_ch_result_Sextans_4__write;
  wire [512:0] fifo_C_ch_result_Sextans_5__dout;
  wire fifo_C_ch_result_Sextans_5__empty_n;
  wire fifo_C_ch_result_Sextans_5__read;
  wire [512:0] fifo_C_ch_result_Sextans_5__din;
  wire fifo_C_ch_result_Sextans_5__full_n;
  wire fifo_C_ch_result_Sextans_5__write;
  wire [512:0] fifo_C_ch_result_Sextans_6__dout;
  wire fifo_C_ch_result_Sextans_6__empty_n;
  wire fifo_C_ch_result_Sextans_6__read;
  wire [512:0] fifo_C_ch_result_Sextans_6__din;
  wire fifo_C_ch_result_Sextans_6__full_n;
  wire fifo_C_ch_result_Sextans_6__write;
  wire [512:0] fifo_C_ch_result_Sextans_7__dout;
  wire fifo_C_ch_result_Sextans_7__empty_n;
  wire fifo_C_ch_result_Sextans_7__read;
  wire [512:0] fifo_C_ch_result_Sextans_7__din;
  wire fifo_C_ch_result_Sextans_7__full_n;
  wire fifo_C_ch_result_Sextans_7__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_0__dout;
  wire fifo_C_ch_result_alpha_Sextans_0__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_0__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_0__din;
  wire fifo_C_ch_result_alpha_Sextans_0__full_n;
  wire fifo_C_ch_result_alpha_Sextans_0__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_1__dout;
  wire fifo_C_ch_result_alpha_Sextans_1__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_1__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_1__din;
  wire fifo_C_ch_result_alpha_Sextans_1__full_n;
  wire fifo_C_ch_result_alpha_Sextans_1__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_2__dout;
  wire fifo_C_ch_result_alpha_Sextans_2__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_2__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_2__din;
  wire fifo_C_ch_result_alpha_Sextans_2__full_n;
  wire fifo_C_ch_result_alpha_Sextans_2__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_3__dout;
  wire fifo_C_ch_result_alpha_Sextans_3__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_3__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_3__din;
  wire fifo_C_ch_result_alpha_Sextans_3__full_n;
  wire fifo_C_ch_result_alpha_Sextans_3__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_4__dout;
  wire fifo_C_ch_result_alpha_Sextans_4__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_4__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_4__din;
  wire fifo_C_ch_result_alpha_Sextans_4__full_n;
  wire fifo_C_ch_result_alpha_Sextans_4__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_5__dout;
  wire fifo_C_ch_result_alpha_Sextans_5__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_5__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_5__din;
  wire fifo_C_ch_result_alpha_Sextans_5__full_n;
  wire fifo_C_ch_result_alpha_Sextans_5__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_6__dout;
  wire fifo_C_ch_result_alpha_Sextans_6__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_6__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_6__din;
  wire fifo_C_ch_result_alpha_Sextans_6__full_n;
  wire fifo_C_ch_result_alpha_Sextans_6__write;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_7__dout;
  wire fifo_C_ch_result_alpha_Sextans_7__empty_n;
  wire fifo_C_ch_result_alpha_Sextans_7__read;
  wire [512:0] fifo_C_ch_result_alpha_Sextans_7__din;
  wire fifo_C_ch_result_alpha_Sextans_7__full_n;
  wire fifo_C_ch_result_alpha_Sextans_7__write;
  wire [256:0] fifo_C_pe_Sextans_0__dout;
  wire fifo_C_pe_Sextans_0__empty_n;
  wire fifo_C_pe_Sextans_0__read;
  wire [256:0] fifo_C_pe_Sextans_0__din;
  wire fifo_C_pe_Sextans_0__full_n;
  wire fifo_C_pe_Sextans_0__write;
  wire [256:0] fifo_C_pe_Sextans_10__dout;
  wire fifo_C_pe_Sextans_10__empty_n;
  wire fifo_C_pe_Sextans_10__read;
  wire [256:0] fifo_C_pe_Sextans_10__din;
  wire fifo_C_pe_Sextans_10__full_n;
  wire fifo_C_pe_Sextans_10__write;
  wire [256:0] fifo_C_pe_Sextans_11__dout;
  wire fifo_C_pe_Sextans_11__empty_n;
  wire fifo_C_pe_Sextans_11__read;
  wire [256:0] fifo_C_pe_Sextans_11__din;
  wire fifo_C_pe_Sextans_11__full_n;
  wire fifo_C_pe_Sextans_11__write;
  wire [256:0] fifo_C_pe_Sextans_12__dout;
  wire fifo_C_pe_Sextans_12__empty_n;
  wire fifo_C_pe_Sextans_12__read;
  wire [256:0] fifo_C_pe_Sextans_12__din;
  wire fifo_C_pe_Sextans_12__full_n;
  wire fifo_C_pe_Sextans_12__write;
  wire [256:0] fifo_C_pe_Sextans_13__dout;
  wire fifo_C_pe_Sextans_13__empty_n;
  wire fifo_C_pe_Sextans_13__read;
  wire [256:0] fifo_C_pe_Sextans_13__din;
  wire fifo_C_pe_Sextans_13__full_n;
  wire fifo_C_pe_Sextans_13__write;
  wire [256:0] fifo_C_pe_Sextans_14__dout;
  wire fifo_C_pe_Sextans_14__empty_n;
  wire fifo_C_pe_Sextans_14__read;
  wire [256:0] fifo_C_pe_Sextans_14__din;
  wire fifo_C_pe_Sextans_14__full_n;
  wire fifo_C_pe_Sextans_14__write;
  wire [256:0] fifo_C_pe_Sextans_15__dout;
  wire fifo_C_pe_Sextans_15__empty_n;
  wire fifo_C_pe_Sextans_15__read;
  wire [256:0] fifo_C_pe_Sextans_15__din;
  wire fifo_C_pe_Sextans_15__full_n;
  wire fifo_C_pe_Sextans_15__write;
  wire [256:0] fifo_C_pe_Sextans_1__dout;
  wire fifo_C_pe_Sextans_1__empty_n;
  wire fifo_C_pe_Sextans_1__read;
  wire [256:0] fifo_C_pe_Sextans_1__din;
  wire fifo_C_pe_Sextans_1__full_n;
  wire fifo_C_pe_Sextans_1__write;
  wire [256:0] fifo_C_pe_Sextans_2__dout;
  wire fifo_C_pe_Sextans_2__empty_n;
  wire fifo_C_pe_Sextans_2__read;
  wire [256:0] fifo_C_pe_Sextans_2__din;
  wire fifo_C_pe_Sextans_2__full_n;
  wire fifo_C_pe_Sextans_2__write;
  wire [256:0] fifo_C_pe_Sextans_3__dout;
  wire fifo_C_pe_Sextans_3__empty_n;
  wire fifo_C_pe_Sextans_3__read;
  wire [256:0] fifo_C_pe_Sextans_3__din;
  wire fifo_C_pe_Sextans_3__full_n;
  wire fifo_C_pe_Sextans_3__write;
  wire [256:0] fifo_C_pe_Sextans_4__dout;
  wire fifo_C_pe_Sextans_4__empty_n;
  wire fifo_C_pe_Sextans_4__read;
  wire [256:0] fifo_C_pe_Sextans_4__din;
  wire fifo_C_pe_Sextans_4__full_n;
  wire fifo_C_pe_Sextans_4__write;
  wire [256:0] fifo_C_pe_Sextans_5__dout;
  wire fifo_C_pe_Sextans_5__empty_n;
  wire fifo_C_pe_Sextans_5__read;
  wire [256:0] fifo_C_pe_Sextans_5__din;
  wire fifo_C_pe_Sextans_5__full_n;
  wire fifo_C_pe_Sextans_5__write;
  wire [256:0] fifo_C_pe_Sextans_6__dout;
  wire fifo_C_pe_Sextans_6__empty_n;
  wire fifo_C_pe_Sextans_6__read;
  wire [256:0] fifo_C_pe_Sextans_6__din;
  wire fifo_C_pe_Sextans_6__full_n;
  wire fifo_C_pe_Sextans_6__write;
  wire [256:0] fifo_C_pe_Sextans_7__dout;
  wire fifo_C_pe_Sextans_7__empty_n;
  wire fifo_C_pe_Sextans_7__read;
  wire [256:0] fifo_C_pe_Sextans_7__din;
  wire fifo_C_pe_Sextans_7__full_n;
  wire fifo_C_pe_Sextans_7__write;
  wire [256:0] fifo_C_pe_Sextans_8__dout;
  wire fifo_C_pe_Sextans_8__empty_n;
  wire fifo_C_pe_Sextans_8__read;
  wire [256:0] fifo_C_pe_Sextans_8__din;
  wire fifo_C_pe_Sextans_8__full_n;
  wire fifo_C_pe_Sextans_8__write;
  wire [256:0] fifo_C_pe_Sextans_9__dout;
  wire fifo_C_pe_Sextans_9__empty_n;
  wire fifo_C_pe_Sextans_9__read;
  wire [256:0] fifo_C_pe_Sextans_9__din;
  wire fifo_C_pe_Sextans_9__full_n;
  wire fifo_C_pe_Sextans_9__write;
  wire [512:0] fifo_C_read_in_Sextans_0__dout;
  wire fifo_C_read_in_Sextans_0__empty_n;
  wire fifo_C_read_in_Sextans_0__read;
  wire [512:0] fifo_C_read_in_Sextans_0__din;
  wire fifo_C_read_in_Sextans_0__full_n;
  wire fifo_C_read_in_Sextans_0__write;
  wire [512:0] fifo_C_read_in_Sextans_1__dout;
  wire fifo_C_read_in_Sextans_1__empty_n;
  wire fifo_C_read_in_Sextans_1__read;
  wire [512:0] fifo_C_read_in_Sextans_1__din;
  wire fifo_C_read_in_Sextans_1__full_n;
  wire fifo_C_read_in_Sextans_1__write;
  wire [512:0] fifo_C_read_in_Sextans_2__dout;
  wire fifo_C_read_in_Sextans_2__empty_n;
  wire fifo_C_read_in_Sextans_2__read;
  wire [512:0] fifo_C_read_in_Sextans_2__din;
  wire fifo_C_read_in_Sextans_2__full_n;
  wire fifo_C_read_in_Sextans_2__write;
  wire [512:0] fifo_C_read_in_Sextans_3__dout;
  wire fifo_C_read_in_Sextans_3__empty_n;
  wire fifo_C_read_in_Sextans_3__read;
  wire [512:0] fifo_C_read_in_Sextans_3__din;
  wire fifo_C_read_in_Sextans_3__full_n;
  wire fifo_C_read_in_Sextans_3__write;
  wire [512:0] fifo_C_read_in_Sextans_4__dout;
  wire fifo_C_read_in_Sextans_4__empty_n;
  wire fifo_C_read_in_Sextans_4__read;
  wire [512:0] fifo_C_read_in_Sextans_4__din;
  wire fifo_C_read_in_Sextans_4__full_n;
  wire fifo_C_read_in_Sextans_4__write;
  wire [512:0] fifo_C_read_in_Sextans_5__dout;
  wire fifo_C_read_in_Sextans_5__empty_n;
  wire fifo_C_read_in_Sextans_5__read;
  wire [512:0] fifo_C_read_in_Sextans_5__din;
  wire fifo_C_read_in_Sextans_5__full_n;
  wire fifo_C_read_in_Sextans_5__write;
  wire [512:0] fifo_C_read_in_Sextans_6__dout;
  wire fifo_C_read_in_Sextans_6__empty_n;
  wire fifo_C_read_in_Sextans_6__read;
  wire [512:0] fifo_C_read_in_Sextans_6__din;
  wire fifo_C_read_in_Sextans_6__full_n;
  wire fifo_C_read_in_Sextans_6__write;
  wire [512:0] fifo_C_read_in_Sextans_7__dout;
  wire fifo_C_read_in_Sextans_7__empty_n;
  wire fifo_C_read_in_Sextans_7__read;
  wire [512:0] fifo_C_read_in_Sextans_7__din;
  wire fifo_C_read_in_Sextans_7__full_n;
  wire fifo_C_read_in_Sextans_7__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_0__dout;
  wire fifo_C_read_in_beta_Sextans_0__empty_n;
  wire fifo_C_read_in_beta_Sextans_0__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_0__din;
  wire fifo_C_read_in_beta_Sextans_0__full_n;
  wire fifo_C_read_in_beta_Sextans_0__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_1__dout;
  wire fifo_C_read_in_beta_Sextans_1__empty_n;
  wire fifo_C_read_in_beta_Sextans_1__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_1__din;
  wire fifo_C_read_in_beta_Sextans_1__full_n;
  wire fifo_C_read_in_beta_Sextans_1__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_2__dout;
  wire fifo_C_read_in_beta_Sextans_2__empty_n;
  wire fifo_C_read_in_beta_Sextans_2__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_2__din;
  wire fifo_C_read_in_beta_Sextans_2__full_n;
  wire fifo_C_read_in_beta_Sextans_2__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_3__dout;
  wire fifo_C_read_in_beta_Sextans_3__empty_n;
  wire fifo_C_read_in_beta_Sextans_3__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_3__din;
  wire fifo_C_read_in_beta_Sextans_3__full_n;
  wire fifo_C_read_in_beta_Sextans_3__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_4__dout;
  wire fifo_C_read_in_beta_Sextans_4__empty_n;
  wire fifo_C_read_in_beta_Sextans_4__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_4__din;
  wire fifo_C_read_in_beta_Sextans_4__full_n;
  wire fifo_C_read_in_beta_Sextans_4__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_5__dout;
  wire fifo_C_read_in_beta_Sextans_5__empty_n;
  wire fifo_C_read_in_beta_Sextans_5__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_5__din;
  wire fifo_C_read_in_beta_Sextans_5__full_n;
  wire fifo_C_read_in_beta_Sextans_5__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_6__dout;
  wire fifo_C_read_in_beta_Sextans_6__empty_n;
  wire fifo_C_read_in_beta_Sextans_6__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_6__din;
  wire fifo_C_read_in_beta_Sextans_6__full_n;
  wire fifo_C_read_in_beta_Sextans_6__write;
  wire [512:0] fifo_C_read_in_beta_Sextans_7__dout;
  wire fifo_C_read_in_beta_Sextans_7__empty_n;
  wire fifo_C_read_in_beta_Sextans_7__read;
  wire [512:0] fifo_C_read_in_beta_Sextans_7__din;
  wire fifo_C_read_in_beta_Sextans_7__full_n;
  wire fifo_C_read_in_beta_Sextans_7__write;
  wire [274:0] fifo_aBvec_Sextans_0__dout;
  wire fifo_aBvec_Sextans_0__empty_n;
  wire fifo_aBvec_Sextans_0__read;
  wire [274:0] fifo_aBvec_Sextans_0__din;
  wire fifo_aBvec_Sextans_0__full_n;
  wire fifo_aBvec_Sextans_0__write;
  wire [274:0] fifo_aBvec_Sextans_10__dout;
  wire fifo_aBvec_Sextans_10__empty_n;
  wire fifo_aBvec_Sextans_10__read;
  wire [274:0] fifo_aBvec_Sextans_10__din;
  wire fifo_aBvec_Sextans_10__full_n;
  wire fifo_aBvec_Sextans_10__write;
  wire [274:0] fifo_aBvec_Sextans_11__dout;
  wire fifo_aBvec_Sextans_11__empty_n;
  wire fifo_aBvec_Sextans_11__read;
  wire [274:0] fifo_aBvec_Sextans_11__din;
  wire fifo_aBvec_Sextans_11__full_n;
  wire fifo_aBvec_Sextans_11__write;
  wire [274:0] fifo_aBvec_Sextans_12__dout;
  wire fifo_aBvec_Sextans_12__empty_n;
  wire fifo_aBvec_Sextans_12__read;
  wire [274:0] fifo_aBvec_Sextans_12__din;
  wire fifo_aBvec_Sextans_12__full_n;
  wire fifo_aBvec_Sextans_12__write;
  wire [274:0] fifo_aBvec_Sextans_13__dout;
  wire fifo_aBvec_Sextans_13__empty_n;
  wire fifo_aBvec_Sextans_13__read;
  wire [274:0] fifo_aBvec_Sextans_13__din;
  wire fifo_aBvec_Sextans_13__full_n;
  wire fifo_aBvec_Sextans_13__write;
  wire [274:0] fifo_aBvec_Sextans_14__dout;
  wire fifo_aBvec_Sextans_14__empty_n;
  wire fifo_aBvec_Sextans_14__read;
  wire [274:0] fifo_aBvec_Sextans_14__din;
  wire fifo_aBvec_Sextans_14__full_n;
  wire fifo_aBvec_Sextans_14__write;
  wire [274:0] fifo_aBvec_Sextans_15__dout;
  wire fifo_aBvec_Sextans_15__empty_n;
  wire fifo_aBvec_Sextans_15__read;
  wire [274:0] fifo_aBvec_Sextans_15__din;
  wire fifo_aBvec_Sextans_15__full_n;
  wire fifo_aBvec_Sextans_15__write;
  wire [274:0] fifo_aBvec_Sextans_16__dout;
  wire fifo_aBvec_Sextans_16__empty_n;
  wire fifo_aBvec_Sextans_16__read;
  wire [274:0] fifo_aBvec_Sextans_16__din;
  wire fifo_aBvec_Sextans_16__full_n;
  wire fifo_aBvec_Sextans_16__write;
  wire [274:0] fifo_aBvec_Sextans_17__dout;
  wire fifo_aBvec_Sextans_17__empty_n;
  wire fifo_aBvec_Sextans_17__read;
  wire [274:0] fifo_aBvec_Sextans_17__din;
  wire fifo_aBvec_Sextans_17__full_n;
  wire fifo_aBvec_Sextans_17__write;
  wire [274:0] fifo_aBvec_Sextans_18__dout;
  wire fifo_aBvec_Sextans_18__empty_n;
  wire fifo_aBvec_Sextans_18__read;
  wire [274:0] fifo_aBvec_Sextans_18__din;
  wire fifo_aBvec_Sextans_18__full_n;
  wire fifo_aBvec_Sextans_18__write;
  wire [274:0] fifo_aBvec_Sextans_19__dout;
  wire fifo_aBvec_Sextans_19__empty_n;
  wire fifo_aBvec_Sextans_19__read;
  wire [274:0] fifo_aBvec_Sextans_19__din;
  wire fifo_aBvec_Sextans_19__full_n;
  wire fifo_aBvec_Sextans_19__write;
  wire [274:0] fifo_aBvec_Sextans_1__dout;
  wire fifo_aBvec_Sextans_1__empty_n;
  wire fifo_aBvec_Sextans_1__read;
  wire [274:0] fifo_aBvec_Sextans_1__din;
  wire fifo_aBvec_Sextans_1__full_n;
  wire fifo_aBvec_Sextans_1__write;
  wire [274:0] fifo_aBvec_Sextans_20__dout;
  wire fifo_aBvec_Sextans_20__empty_n;
  wire fifo_aBvec_Sextans_20__read;
  wire [274:0] fifo_aBvec_Sextans_20__din;
  wire fifo_aBvec_Sextans_20__full_n;
  wire fifo_aBvec_Sextans_20__write;
  wire [274:0] fifo_aBvec_Sextans_21__dout;
  wire fifo_aBvec_Sextans_21__empty_n;
  wire fifo_aBvec_Sextans_21__read;
  wire [274:0] fifo_aBvec_Sextans_21__din;
  wire fifo_aBvec_Sextans_21__full_n;
  wire fifo_aBvec_Sextans_21__write;
  wire [274:0] fifo_aBvec_Sextans_22__dout;
  wire fifo_aBvec_Sextans_22__empty_n;
  wire fifo_aBvec_Sextans_22__read;
  wire [274:0] fifo_aBvec_Sextans_22__din;
  wire fifo_aBvec_Sextans_22__full_n;
  wire fifo_aBvec_Sextans_22__write;
  wire [274:0] fifo_aBvec_Sextans_23__dout;
  wire fifo_aBvec_Sextans_23__empty_n;
  wire fifo_aBvec_Sextans_23__read;
  wire [274:0] fifo_aBvec_Sextans_23__din;
  wire fifo_aBvec_Sextans_23__full_n;
  wire fifo_aBvec_Sextans_23__write;
  wire [274:0] fifo_aBvec_Sextans_24__dout;
  wire fifo_aBvec_Sextans_24__empty_n;
  wire fifo_aBvec_Sextans_24__read;
  wire [274:0] fifo_aBvec_Sextans_24__din;
  wire fifo_aBvec_Sextans_24__full_n;
  wire fifo_aBvec_Sextans_24__write;
  wire [274:0] fifo_aBvec_Sextans_25__dout;
  wire fifo_aBvec_Sextans_25__empty_n;
  wire fifo_aBvec_Sextans_25__read;
  wire [274:0] fifo_aBvec_Sextans_25__din;
  wire fifo_aBvec_Sextans_25__full_n;
  wire fifo_aBvec_Sextans_25__write;
  wire [274:0] fifo_aBvec_Sextans_26__dout;
  wire fifo_aBvec_Sextans_26__empty_n;
  wire fifo_aBvec_Sextans_26__read;
  wire [274:0] fifo_aBvec_Sextans_26__din;
  wire fifo_aBvec_Sextans_26__full_n;
  wire fifo_aBvec_Sextans_26__write;
  wire [274:0] fifo_aBvec_Sextans_27__dout;
  wire fifo_aBvec_Sextans_27__empty_n;
  wire fifo_aBvec_Sextans_27__read;
  wire [274:0] fifo_aBvec_Sextans_27__din;
  wire fifo_aBvec_Sextans_27__full_n;
  wire fifo_aBvec_Sextans_27__write;
  wire [274:0] fifo_aBvec_Sextans_28__dout;
  wire fifo_aBvec_Sextans_28__empty_n;
  wire fifo_aBvec_Sextans_28__read;
  wire [274:0] fifo_aBvec_Sextans_28__din;
  wire fifo_aBvec_Sextans_28__full_n;
  wire fifo_aBvec_Sextans_28__write;
  wire [274:0] fifo_aBvec_Sextans_29__dout;
  wire fifo_aBvec_Sextans_29__empty_n;
  wire fifo_aBvec_Sextans_29__read;
  wire [274:0] fifo_aBvec_Sextans_29__din;
  wire fifo_aBvec_Sextans_29__full_n;
  wire fifo_aBvec_Sextans_29__write;
  wire [274:0] fifo_aBvec_Sextans_2__dout;
  wire fifo_aBvec_Sextans_2__empty_n;
  wire fifo_aBvec_Sextans_2__read;
  wire [274:0] fifo_aBvec_Sextans_2__din;
  wire fifo_aBvec_Sextans_2__full_n;
  wire fifo_aBvec_Sextans_2__write;
  wire [274:0] fifo_aBvec_Sextans_30__dout;
  wire fifo_aBvec_Sextans_30__empty_n;
  wire fifo_aBvec_Sextans_30__read;
  wire [274:0] fifo_aBvec_Sextans_30__din;
  wire fifo_aBvec_Sextans_30__full_n;
  wire fifo_aBvec_Sextans_30__write;
  wire [274:0] fifo_aBvec_Sextans_31__dout;
  wire fifo_aBvec_Sextans_31__empty_n;
  wire fifo_aBvec_Sextans_31__read;
  wire [274:0] fifo_aBvec_Sextans_31__din;
  wire fifo_aBvec_Sextans_31__full_n;
  wire fifo_aBvec_Sextans_31__write;
  wire [274:0] fifo_aBvec_Sextans_32__dout;
  wire fifo_aBvec_Sextans_32__empty_n;
  wire fifo_aBvec_Sextans_32__read;
  wire [274:0] fifo_aBvec_Sextans_32__din;
  wire fifo_aBvec_Sextans_32__full_n;
  wire fifo_aBvec_Sextans_32__write;
  wire [274:0] fifo_aBvec_Sextans_33__dout;
  wire fifo_aBvec_Sextans_33__empty_n;
  wire fifo_aBvec_Sextans_33__read;
  wire [274:0] fifo_aBvec_Sextans_33__din;
  wire fifo_aBvec_Sextans_33__full_n;
  wire fifo_aBvec_Sextans_33__write;
  wire [274:0] fifo_aBvec_Sextans_34__dout;
  wire fifo_aBvec_Sextans_34__empty_n;
  wire fifo_aBvec_Sextans_34__read;
  wire [274:0] fifo_aBvec_Sextans_34__din;
  wire fifo_aBvec_Sextans_34__full_n;
  wire fifo_aBvec_Sextans_34__write;
  wire [274:0] fifo_aBvec_Sextans_35__dout;
  wire fifo_aBvec_Sextans_35__empty_n;
  wire fifo_aBvec_Sextans_35__read;
  wire [274:0] fifo_aBvec_Sextans_35__din;
  wire fifo_aBvec_Sextans_35__full_n;
  wire fifo_aBvec_Sextans_35__write;
  wire [274:0] fifo_aBvec_Sextans_36__dout;
  wire fifo_aBvec_Sextans_36__empty_n;
  wire fifo_aBvec_Sextans_36__read;
  wire [274:0] fifo_aBvec_Sextans_36__din;
  wire fifo_aBvec_Sextans_36__full_n;
  wire fifo_aBvec_Sextans_36__write;
  wire [274:0] fifo_aBvec_Sextans_37__dout;
  wire fifo_aBvec_Sextans_37__empty_n;
  wire fifo_aBvec_Sextans_37__read;
  wire [274:0] fifo_aBvec_Sextans_37__din;
  wire fifo_aBvec_Sextans_37__full_n;
  wire fifo_aBvec_Sextans_37__write;
  wire [274:0] fifo_aBvec_Sextans_38__dout;
  wire fifo_aBvec_Sextans_38__empty_n;
  wire fifo_aBvec_Sextans_38__read;
  wire [274:0] fifo_aBvec_Sextans_38__din;
  wire fifo_aBvec_Sextans_38__full_n;
  wire fifo_aBvec_Sextans_38__write;
  wire [274:0] fifo_aBvec_Sextans_39__dout;
  wire fifo_aBvec_Sextans_39__empty_n;
  wire fifo_aBvec_Sextans_39__read;
  wire [274:0] fifo_aBvec_Sextans_39__din;
  wire fifo_aBvec_Sextans_39__full_n;
  wire fifo_aBvec_Sextans_39__write;
  wire [274:0] fifo_aBvec_Sextans_3__dout;
  wire fifo_aBvec_Sextans_3__empty_n;
  wire fifo_aBvec_Sextans_3__read;
  wire [274:0] fifo_aBvec_Sextans_3__din;
  wire fifo_aBvec_Sextans_3__full_n;
  wire fifo_aBvec_Sextans_3__write;
  wire [274:0] fifo_aBvec_Sextans_40__dout;
  wire fifo_aBvec_Sextans_40__empty_n;
  wire fifo_aBvec_Sextans_40__read;
  wire [274:0] fifo_aBvec_Sextans_40__din;
  wire fifo_aBvec_Sextans_40__full_n;
  wire fifo_aBvec_Sextans_40__write;
  wire [274:0] fifo_aBvec_Sextans_41__dout;
  wire fifo_aBvec_Sextans_41__empty_n;
  wire fifo_aBvec_Sextans_41__read;
  wire [274:0] fifo_aBvec_Sextans_41__din;
  wire fifo_aBvec_Sextans_41__full_n;
  wire fifo_aBvec_Sextans_41__write;
  wire [274:0] fifo_aBvec_Sextans_42__dout;
  wire fifo_aBvec_Sextans_42__empty_n;
  wire fifo_aBvec_Sextans_42__read;
  wire [274:0] fifo_aBvec_Sextans_42__din;
  wire fifo_aBvec_Sextans_42__full_n;
  wire fifo_aBvec_Sextans_42__write;
  wire [274:0] fifo_aBvec_Sextans_43__dout;
  wire fifo_aBvec_Sextans_43__empty_n;
  wire fifo_aBvec_Sextans_43__read;
  wire [274:0] fifo_aBvec_Sextans_43__din;
  wire fifo_aBvec_Sextans_43__full_n;
  wire fifo_aBvec_Sextans_43__write;
  wire [274:0] fifo_aBvec_Sextans_44__dout;
  wire fifo_aBvec_Sextans_44__empty_n;
  wire fifo_aBvec_Sextans_44__read;
  wire [274:0] fifo_aBvec_Sextans_44__din;
  wire fifo_aBvec_Sextans_44__full_n;
  wire fifo_aBvec_Sextans_44__write;
  wire [274:0] fifo_aBvec_Sextans_45__dout;
  wire fifo_aBvec_Sextans_45__empty_n;
  wire fifo_aBvec_Sextans_45__read;
  wire [274:0] fifo_aBvec_Sextans_45__din;
  wire fifo_aBvec_Sextans_45__full_n;
  wire fifo_aBvec_Sextans_45__write;
  wire [274:0] fifo_aBvec_Sextans_46__dout;
  wire fifo_aBvec_Sextans_46__empty_n;
  wire fifo_aBvec_Sextans_46__read;
  wire [274:0] fifo_aBvec_Sextans_46__din;
  wire fifo_aBvec_Sextans_46__full_n;
  wire fifo_aBvec_Sextans_46__write;
  wire [274:0] fifo_aBvec_Sextans_47__dout;
  wire fifo_aBvec_Sextans_47__empty_n;
  wire fifo_aBvec_Sextans_47__read;
  wire [274:0] fifo_aBvec_Sextans_47__din;
  wire fifo_aBvec_Sextans_47__full_n;
  wire fifo_aBvec_Sextans_47__write;
  wire [274:0] fifo_aBvec_Sextans_48__dout;
  wire fifo_aBvec_Sextans_48__empty_n;
  wire fifo_aBvec_Sextans_48__read;
  wire [274:0] fifo_aBvec_Sextans_48__din;
  wire fifo_aBvec_Sextans_48__full_n;
  wire fifo_aBvec_Sextans_48__write;
  wire [274:0] fifo_aBvec_Sextans_49__dout;
  wire fifo_aBvec_Sextans_49__empty_n;
  wire fifo_aBvec_Sextans_49__read;
  wire [274:0] fifo_aBvec_Sextans_49__din;
  wire fifo_aBvec_Sextans_49__full_n;
  wire fifo_aBvec_Sextans_49__write;
  wire [274:0] fifo_aBvec_Sextans_4__dout;
  wire fifo_aBvec_Sextans_4__empty_n;
  wire fifo_aBvec_Sextans_4__read;
  wire [274:0] fifo_aBvec_Sextans_4__din;
  wire fifo_aBvec_Sextans_4__full_n;
  wire fifo_aBvec_Sextans_4__write;
  wire [274:0] fifo_aBvec_Sextans_50__dout;
  wire fifo_aBvec_Sextans_50__empty_n;
  wire fifo_aBvec_Sextans_50__read;
  wire [274:0] fifo_aBvec_Sextans_50__din;
  wire fifo_aBvec_Sextans_50__full_n;
  wire fifo_aBvec_Sextans_50__write;
  wire [274:0] fifo_aBvec_Sextans_51__dout;
  wire fifo_aBvec_Sextans_51__empty_n;
  wire fifo_aBvec_Sextans_51__read;
  wire [274:0] fifo_aBvec_Sextans_51__din;
  wire fifo_aBvec_Sextans_51__full_n;
  wire fifo_aBvec_Sextans_51__write;
  wire [274:0] fifo_aBvec_Sextans_52__dout;
  wire fifo_aBvec_Sextans_52__empty_n;
  wire fifo_aBvec_Sextans_52__read;
  wire [274:0] fifo_aBvec_Sextans_52__din;
  wire fifo_aBvec_Sextans_52__full_n;
  wire fifo_aBvec_Sextans_52__write;
  wire [274:0] fifo_aBvec_Sextans_53__dout;
  wire fifo_aBvec_Sextans_53__empty_n;
  wire fifo_aBvec_Sextans_53__read;
  wire [274:0] fifo_aBvec_Sextans_53__din;
  wire fifo_aBvec_Sextans_53__full_n;
  wire fifo_aBvec_Sextans_53__write;
  wire [274:0] fifo_aBvec_Sextans_54__dout;
  wire fifo_aBvec_Sextans_54__empty_n;
  wire fifo_aBvec_Sextans_54__read;
  wire [274:0] fifo_aBvec_Sextans_54__din;
  wire fifo_aBvec_Sextans_54__full_n;
  wire fifo_aBvec_Sextans_54__write;
  wire [274:0] fifo_aBvec_Sextans_55__dout;
  wire fifo_aBvec_Sextans_55__empty_n;
  wire fifo_aBvec_Sextans_55__read;
  wire [274:0] fifo_aBvec_Sextans_55__din;
  wire fifo_aBvec_Sextans_55__full_n;
  wire fifo_aBvec_Sextans_55__write;
  wire [274:0] fifo_aBvec_Sextans_56__dout;
  wire fifo_aBvec_Sextans_56__empty_n;
  wire fifo_aBvec_Sextans_56__read;
  wire [274:0] fifo_aBvec_Sextans_56__din;
  wire fifo_aBvec_Sextans_56__full_n;
  wire fifo_aBvec_Sextans_56__write;
  wire [274:0] fifo_aBvec_Sextans_57__dout;
  wire fifo_aBvec_Sextans_57__empty_n;
  wire fifo_aBvec_Sextans_57__read;
  wire [274:0] fifo_aBvec_Sextans_57__din;
  wire fifo_aBvec_Sextans_57__full_n;
  wire fifo_aBvec_Sextans_57__write;
  wire [274:0] fifo_aBvec_Sextans_58__dout;
  wire fifo_aBvec_Sextans_58__empty_n;
  wire fifo_aBvec_Sextans_58__read;
  wire [274:0] fifo_aBvec_Sextans_58__din;
  wire fifo_aBvec_Sextans_58__full_n;
  wire fifo_aBvec_Sextans_58__write;
  wire [274:0] fifo_aBvec_Sextans_59__dout;
  wire fifo_aBvec_Sextans_59__empty_n;
  wire fifo_aBvec_Sextans_59__read;
  wire [274:0] fifo_aBvec_Sextans_59__din;
  wire fifo_aBvec_Sextans_59__full_n;
  wire fifo_aBvec_Sextans_59__write;
  wire [274:0] fifo_aBvec_Sextans_5__dout;
  wire fifo_aBvec_Sextans_5__empty_n;
  wire fifo_aBvec_Sextans_5__read;
  wire [274:0] fifo_aBvec_Sextans_5__din;
  wire fifo_aBvec_Sextans_5__full_n;
  wire fifo_aBvec_Sextans_5__write;
  wire [274:0] fifo_aBvec_Sextans_60__dout;
  wire fifo_aBvec_Sextans_60__empty_n;
  wire fifo_aBvec_Sextans_60__read;
  wire [274:0] fifo_aBvec_Sextans_60__din;
  wire fifo_aBvec_Sextans_60__full_n;
  wire fifo_aBvec_Sextans_60__write;
  wire [274:0] fifo_aBvec_Sextans_61__dout;
  wire fifo_aBvec_Sextans_61__empty_n;
  wire fifo_aBvec_Sextans_61__read;
  wire [274:0] fifo_aBvec_Sextans_61__din;
  wire fifo_aBvec_Sextans_61__full_n;
  wire fifo_aBvec_Sextans_61__write;
  wire [274:0] fifo_aBvec_Sextans_62__dout;
  wire fifo_aBvec_Sextans_62__empty_n;
  wire fifo_aBvec_Sextans_62__read;
  wire [274:0] fifo_aBvec_Sextans_62__din;
  wire fifo_aBvec_Sextans_62__full_n;
  wire fifo_aBvec_Sextans_62__write;
  wire [274:0] fifo_aBvec_Sextans_63__dout;
  wire fifo_aBvec_Sextans_63__empty_n;
  wire fifo_aBvec_Sextans_63__read;
  wire [274:0] fifo_aBvec_Sextans_63__din;
  wire fifo_aBvec_Sextans_63__full_n;
  wire fifo_aBvec_Sextans_63__write;
  wire [274:0] fifo_aBvec_Sextans_6__dout;
  wire fifo_aBvec_Sextans_6__empty_n;
  wire fifo_aBvec_Sextans_6__read;
  wire [274:0] fifo_aBvec_Sextans_6__din;
  wire fifo_aBvec_Sextans_6__full_n;
  wire fifo_aBvec_Sextans_6__write;
  wire [274:0] fifo_aBvec_Sextans_7__dout;
  wire fifo_aBvec_Sextans_7__empty_n;
  wire fifo_aBvec_Sextans_7__read;
  wire [274:0] fifo_aBvec_Sextans_7__din;
  wire fifo_aBvec_Sextans_7__full_n;
  wire fifo_aBvec_Sextans_7__write;
  wire [274:0] fifo_aBvec_Sextans_8__dout;
  wire fifo_aBvec_Sextans_8__empty_n;
  wire fifo_aBvec_Sextans_8__read;
  wire [274:0] fifo_aBvec_Sextans_8__din;
  wire fifo_aBvec_Sextans_8__full_n;
  wire fifo_aBvec_Sextans_8__write;
  wire [274:0] fifo_aBvec_Sextans_9__dout;
  wire fifo_aBvec_Sextans_9__empty_n;
  wire fifo_aBvec_Sextans_9__read;
  wire [274:0] fifo_aBvec_Sextans_9__din;
  wire fifo_aBvec_Sextans_9__full_n;
  wire fifo_aBvec_Sextans_9__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_0__dout;
  wire fifo_edge_list_ptr_Sextans_0__empty_n;
  wire fifo_edge_list_ptr_Sextans_0__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_0__din;
  wire fifo_edge_list_ptr_Sextans_0__full_n;
  wire fifo_edge_list_ptr_Sextans_0__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_10__dout;
  wire fifo_edge_list_ptr_Sextans_10__empty_n;
  wire fifo_edge_list_ptr_Sextans_10__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_10__din;
  wire fifo_edge_list_ptr_Sextans_10__full_n;
  wire fifo_edge_list_ptr_Sextans_10__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_11__dout;
  wire fifo_edge_list_ptr_Sextans_11__empty_n;
  wire fifo_edge_list_ptr_Sextans_11__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_11__din;
  wire fifo_edge_list_ptr_Sextans_11__full_n;
  wire fifo_edge_list_ptr_Sextans_11__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_12__dout;
  wire fifo_edge_list_ptr_Sextans_12__empty_n;
  wire fifo_edge_list_ptr_Sextans_12__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_12__din;
  wire fifo_edge_list_ptr_Sextans_12__full_n;
  wire fifo_edge_list_ptr_Sextans_12__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_13__dout;
  wire fifo_edge_list_ptr_Sextans_13__empty_n;
  wire fifo_edge_list_ptr_Sextans_13__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_13__din;
  wire fifo_edge_list_ptr_Sextans_13__full_n;
  wire fifo_edge_list_ptr_Sextans_13__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_14__dout;
  wire fifo_edge_list_ptr_Sextans_14__empty_n;
  wire fifo_edge_list_ptr_Sextans_14__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_14__din;
  wire fifo_edge_list_ptr_Sextans_14__full_n;
  wire fifo_edge_list_ptr_Sextans_14__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_15__dout;
  wire fifo_edge_list_ptr_Sextans_15__empty_n;
  wire fifo_edge_list_ptr_Sextans_15__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_15__din;
  wire fifo_edge_list_ptr_Sextans_15__full_n;
  wire fifo_edge_list_ptr_Sextans_15__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_16__dout;
  wire fifo_edge_list_ptr_Sextans_16__empty_n;
  wire fifo_edge_list_ptr_Sextans_16__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_16__din;
  wire fifo_edge_list_ptr_Sextans_16__full_n;
  wire fifo_edge_list_ptr_Sextans_16__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_1__dout;
  wire fifo_edge_list_ptr_Sextans_1__empty_n;
  wire fifo_edge_list_ptr_Sextans_1__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_1__din;
  wire fifo_edge_list_ptr_Sextans_1__full_n;
  wire fifo_edge_list_ptr_Sextans_1__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_2__dout;
  wire fifo_edge_list_ptr_Sextans_2__empty_n;
  wire fifo_edge_list_ptr_Sextans_2__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_2__din;
  wire fifo_edge_list_ptr_Sextans_2__full_n;
  wire fifo_edge_list_ptr_Sextans_2__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_3__dout;
  wire fifo_edge_list_ptr_Sextans_3__empty_n;
  wire fifo_edge_list_ptr_Sextans_3__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_3__din;
  wire fifo_edge_list_ptr_Sextans_3__full_n;
  wire fifo_edge_list_ptr_Sextans_3__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_4__dout;
  wire fifo_edge_list_ptr_Sextans_4__empty_n;
  wire fifo_edge_list_ptr_Sextans_4__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_4__din;
  wire fifo_edge_list_ptr_Sextans_4__full_n;
  wire fifo_edge_list_ptr_Sextans_4__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_5__dout;
  wire fifo_edge_list_ptr_Sextans_5__empty_n;
  wire fifo_edge_list_ptr_Sextans_5__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_5__din;
  wire fifo_edge_list_ptr_Sextans_5__full_n;
  wire fifo_edge_list_ptr_Sextans_5__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_6__dout;
  wire fifo_edge_list_ptr_Sextans_6__empty_n;
  wire fifo_edge_list_ptr_Sextans_6__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_6__din;
  wire fifo_edge_list_ptr_Sextans_6__full_n;
  wire fifo_edge_list_ptr_Sextans_6__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_7__dout;
  wire fifo_edge_list_ptr_Sextans_7__empty_n;
  wire fifo_edge_list_ptr_Sextans_7__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_7__din;
  wire fifo_edge_list_ptr_Sextans_7__full_n;
  wire fifo_edge_list_ptr_Sextans_7__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_8__dout;
  wire fifo_edge_list_ptr_Sextans_8__empty_n;
  wire fifo_edge_list_ptr_Sextans_8__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_8__din;
  wire fifo_edge_list_ptr_Sextans_8__full_n;
  wire fifo_edge_list_ptr_Sextans_8__write;
  wire [32:0] fifo_edge_list_ptr_Sextans_9__dout;
  wire fifo_edge_list_ptr_Sextans_9__empty_n;
  wire fifo_edge_list_ptr_Sextans_9__read;
  wire [32:0] fifo_edge_list_ptr_Sextans_9__din;
  wire fifo_edge_list_ptr_Sextans_9__full_n;
  wire fifo_edge_list_ptr_Sextans_9__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_0__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_0__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_0__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_0__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_0__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_0__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_10__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_10__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_10__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_10__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_10__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_10__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_11__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_11__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_11__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_11__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_11__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_11__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_12__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_12__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_12__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_12__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_12__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_12__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_13__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_13__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_13__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_13__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_13__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_13__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_14__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_14__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_14__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_14__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_14__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_14__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_15__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_15__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_15__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_15__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_15__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_15__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_1__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_1__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_1__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_1__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_1__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_1__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_2__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_2__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_2__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_2__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_2__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_2__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_3__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_3__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_3__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_3__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_3__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_3__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_4__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_4__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_4__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_4__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_4__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_4__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_5__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_5__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_5__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_5__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_5__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_5__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_6__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_6__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_6__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_6__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_6__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_6__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_7__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_7__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_7__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_7__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_7__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_7__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_8__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_8__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_8__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_8__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_8__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_8__write;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_9__dout;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_9__empty_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_9__read;
  wire [32:0] fifo_edge_list_ptr_to_Cmtx_Sextans_9__din;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_9__full_n;
  wire fifo_edge_list_ptr_to_Cmtx_Sextans_9__write;
  wire [32:0] wrC_inst_Sextans_0__dout;
  wire wrC_inst_Sextans_0__empty_n;
  wire wrC_inst_Sextans_0__read;
  wire [32:0] wrC_inst_Sextans_0__din;
  wire wrC_inst_Sextans_0__full_n;
  wire wrC_inst_Sextans_0__write;
  wire [32:0] wrC_inst_Sextans_1__dout;
  wire wrC_inst_Sextans_1__empty_n;
  wire wrC_inst_Sextans_1__read;
  wire [32:0] wrC_inst_Sextans_1__din;
  wire wrC_inst_Sextans_1__full_n;
  wire wrC_inst_Sextans_1__write;
  wire [32:0] wrC_inst_Sextans_2__dout;
  wire wrC_inst_Sextans_2__empty_n;
  wire wrC_inst_Sextans_2__read;
  wire [32:0] wrC_inst_Sextans_2__din;
  wire wrC_inst_Sextans_2__full_n;
  wire wrC_inst_Sextans_2__write;
  wire [32:0] wrC_inst_Sextans_3__dout;
  wire wrC_inst_Sextans_3__empty_n;
  wire wrC_inst_Sextans_3__read;
  wire [32:0] wrC_inst_Sextans_3__din;
  wire wrC_inst_Sextans_3__full_n;
  wire wrC_inst_Sextans_3__write;
  wire [32:0] wrC_inst_Sextans_4__dout;
  wire wrC_inst_Sextans_4__empty_n;
  wire wrC_inst_Sextans_4__read;
  wire [32:0] wrC_inst_Sextans_4__din;
  wire wrC_inst_Sextans_4__full_n;
  wire wrC_inst_Sextans_4__write;
  wire [32:0] wrC_inst_Sextans_5__dout;
  wire wrC_inst_Sextans_5__empty_n;
  wire wrC_inst_Sextans_5__read;
  wire [32:0] wrC_inst_Sextans_5__din;
  wire wrC_inst_Sextans_5__full_n;
  wire wrC_inst_Sextans_5__write;
  wire [32:0] wrC_inst_Sextans_6__dout;
  wire wrC_inst_Sextans_6__empty_n;
  wire wrC_inst_Sextans_6__read;
  wire [32:0] wrC_inst_Sextans_6__din;
  wire wrC_inst_Sextans_6__full_n;
  wire wrC_inst_Sextans_6__write;
  wire [32:0] wrC_inst_Sextans_7__dout;
  wire wrC_inst_Sextans_7__empty_n;
  wire wrC_inst_Sextans_7__read;
  wire [32:0] wrC_inst_Sextans_7__din;
  wire wrC_inst_Sextans_7__full_n;
  wire wrC_inst_Sextans_7__write;
  wire FloatvAddFloatv_0__ap_start;
  wire FloatvAddFloatv_1__ap_start;
  wire FloatvAddFloatv_2__ap_start;
  wire FloatvAddFloatv_3__ap_start;
  wire FloatvAddFloatv_4__ap_start;
  wire FloatvAddFloatv_5__ap_start;
  wire FloatvAddFloatv_6__ap_start;
  wire FloatvAddFloatv_7__ap_start;
  wire [31:0] FloatvMultConst_0___M__q0;
  wire [31:0] FloatvMultConst_0___P_N__q0;
  wire [31:0] FloatvMultConst_0___beta_u__q0;
  wire FloatvMultConst_0__ap_start;
  wire FloatvMultConst_0__ap_ready;
  wire FloatvMultConst_0__ap_done;
  wire FloatvMultConst_0__ap_idle;
  wire [31:0] FloatvMultConst_1___M__q0;
  wire [31:0] FloatvMultConst_1___P_N__q0;
  wire [31:0] FloatvMultConst_1___beta_u__q0;
  wire FloatvMultConst_1__ap_start;
  wire FloatvMultConst_1__ap_ready;
  wire FloatvMultConst_1__ap_done;
  wire FloatvMultConst_1__ap_idle;
  wire [31:0] FloatvMultConst_2___M__q0;
  wire [31:0] FloatvMultConst_2___P_N__q0;
  wire [31:0] FloatvMultConst_2___beta_u__q0;
  wire FloatvMultConst_2__ap_start;
  wire FloatvMultConst_2__ap_ready;
  wire FloatvMultConst_2__ap_done;
  wire FloatvMultConst_2__ap_idle;
  wire [31:0] FloatvMultConst_3___M__q0;
  wire [31:0] FloatvMultConst_3___P_N__q0;
  wire [31:0] FloatvMultConst_3___beta_u__q0;
  wire FloatvMultConst_3__ap_start;
  wire FloatvMultConst_3__ap_ready;
  wire FloatvMultConst_3__ap_done;
  wire FloatvMultConst_3__ap_idle;
  wire [31:0] FloatvMultConst_4___M__q0;
  wire [31:0] FloatvMultConst_4___P_N__q0;
  wire [31:0] FloatvMultConst_4___beta_u__q0;
  wire FloatvMultConst_4__ap_start;
  wire FloatvMultConst_4__ap_ready;
  wire FloatvMultConst_4__ap_done;
  wire FloatvMultConst_4__ap_idle;
  wire [31:0] FloatvMultConst_5___M__q0;
  wire [31:0] FloatvMultConst_5___P_N__q0;
  wire [31:0] FloatvMultConst_5___beta_u__q0;
  wire FloatvMultConst_5__ap_start;
  wire FloatvMultConst_5__ap_ready;
  wire FloatvMultConst_5__ap_done;
  wire FloatvMultConst_5__ap_idle;
  wire [31:0] FloatvMultConst_6___M__q0;
  wire [31:0] FloatvMultConst_6___P_N__q0;
  wire [31:0] FloatvMultConst_6___beta_u__q0;
  wire FloatvMultConst_6__ap_start;
  wire FloatvMultConst_6__ap_ready;
  wire FloatvMultConst_6__ap_done;
  wire FloatvMultConst_6__ap_idle;
  wire [31:0] FloatvMultConst_7___M__q0;
  wire [31:0] FloatvMultConst_7___P_N__q0;
  wire [31:0] FloatvMultConst_7___beta_u__q0;
  wire FloatvMultConst_7__ap_start;
  wire FloatvMultConst_7__ap_ready;
  wire FloatvMultConst_7__ap_done;
  wire FloatvMultConst_7__ap_idle;
  wire [31:0] FloatvMultConst_8___M__q0;
  wire [31:0] FloatvMultConst_8___P_N__q0;
  wire [31:0] FloatvMultConst_8___alpha_u__q0;
  wire FloatvMultConst_8__ap_start;
  wire FloatvMultConst_8__ap_ready;
  wire FloatvMultConst_8__ap_done;
  wire FloatvMultConst_8__ap_idle;
  wire [31:0] FloatvMultConst_9___M__q0;
  wire [31:0] FloatvMultConst_9___P_N__q0;
  wire [31:0] FloatvMultConst_9___alpha_u__q0;
  wire FloatvMultConst_9__ap_start;
  wire FloatvMultConst_9__ap_ready;
  wire FloatvMultConst_9__ap_done;
  wire FloatvMultConst_9__ap_idle;
  wire [31:0] FloatvMultConst_10___M__q0;
  wire [31:0] FloatvMultConst_10___P_N__q0;
  wire [31:0] FloatvMultConst_10___alpha_u__q0;
  wire FloatvMultConst_10__ap_start;
  wire FloatvMultConst_10__ap_ready;
  wire FloatvMultConst_10__ap_done;
  wire FloatvMultConst_10__ap_idle;
  wire [31:0] FloatvMultConst_11___M__q0;
  wire [31:0] FloatvMultConst_11___P_N__q0;
  wire [31:0] FloatvMultConst_11___alpha_u__q0;
  wire FloatvMultConst_11__ap_start;
  wire FloatvMultConst_11__ap_ready;
  wire FloatvMultConst_11__ap_done;
  wire FloatvMultConst_11__ap_idle;
  wire [31:0] FloatvMultConst_12___M__q0;
  wire [31:0] FloatvMultConst_12___P_N__q0;
  wire [31:0] FloatvMultConst_12___alpha_u__q0;
  wire FloatvMultConst_12__ap_start;
  wire FloatvMultConst_12__ap_ready;
  wire FloatvMultConst_12__ap_done;
  wire FloatvMultConst_12__ap_idle;
  wire [31:0] FloatvMultConst_13___M__q0;
  wire [31:0] FloatvMultConst_13___P_N__q0;
  wire [31:0] FloatvMultConst_13___alpha_u__q0;
  wire FloatvMultConst_13__ap_start;
  wire FloatvMultConst_13__ap_ready;
  wire FloatvMultConst_13__ap_done;
  wire FloatvMultConst_13__ap_idle;
  wire [31:0] FloatvMultConst_14___M__q0;
  wire [31:0] FloatvMultConst_14___P_N__q0;
  wire [31:0] FloatvMultConst_14___alpha_u__q0;
  wire FloatvMultConst_14__ap_start;
  wire FloatvMultConst_14__ap_ready;
  wire FloatvMultConst_14__ap_done;
  wire FloatvMultConst_14__ap_idle;
  wire [31:0] FloatvMultConst_15___M__q0;
  wire [31:0] FloatvMultConst_15___P_N__q0;
  wire [31:0] FloatvMultConst_15___alpha_u__q0;
  wire FloatvMultConst_15__ap_start;
  wire FloatvMultConst_15__ap_ready;
  wire FloatvMultConst_15__ap_done;
  wire FloatvMultConst_15__ap_idle;
  wire Merger_0__ap_start;
  wire Merger_1__ap_start;
  wire Merger_2__ap_start;
  wire Merger_3__ap_start;
  wire Merger_4__ap_start;
  wire Merger_5__ap_start;
  wire Merger_6__ap_start;
  wire Merger_7__ap_start;
  wire PEG_Bmtx_0__ap_start;
  wire PEG_Bmtx_0__ap_ready;
  wire PEG_Bmtx_0__ap_done;
  wire PEG_Bmtx_0__ap_idle;
  wire PEG_Bmtx_1__ap_start;
  wire PEG_Bmtx_1__ap_ready;
  wire PEG_Bmtx_1__ap_done;
  wire PEG_Bmtx_1__ap_idle;
  wire PEG_Bmtx_2__ap_start;
  wire PEG_Bmtx_2__ap_ready;
  wire PEG_Bmtx_2__ap_done;
  wire PEG_Bmtx_2__ap_idle;
  wire PEG_Bmtx_3__ap_start;
  wire PEG_Bmtx_3__ap_ready;
  wire PEG_Bmtx_3__ap_done;
  wire PEG_Bmtx_3__ap_idle;
  wire PEG_Bmtx_4__ap_start;
  wire PEG_Bmtx_4__ap_ready;
  wire PEG_Bmtx_4__ap_done;
  wire PEG_Bmtx_4__ap_idle;
  wire PEG_Bmtx_5__ap_start;
  wire PEG_Bmtx_5__ap_ready;
  wire PEG_Bmtx_5__ap_done;
  wire PEG_Bmtx_5__ap_idle;
  wire PEG_Bmtx_6__ap_start;
  wire PEG_Bmtx_6__ap_ready;
  wire PEG_Bmtx_6__ap_done;
  wire PEG_Bmtx_6__ap_idle;
  wire PEG_Bmtx_7__ap_start;
  wire PEG_Bmtx_7__ap_ready;
  wire PEG_Bmtx_7__ap_done;
  wire PEG_Bmtx_7__ap_idle;
  wire PEG_Bmtx_8__ap_start;
  wire PEG_Bmtx_8__ap_ready;
  wire PEG_Bmtx_8__ap_done;
  wire PEG_Bmtx_8__ap_idle;
  wire PEG_Bmtx_9__ap_start;
  wire PEG_Bmtx_9__ap_ready;
  wire PEG_Bmtx_9__ap_done;
  wire PEG_Bmtx_9__ap_idle;
  wire PEG_Bmtx_10__ap_start;
  wire PEG_Bmtx_10__ap_ready;
  wire PEG_Bmtx_10__ap_done;
  wire PEG_Bmtx_10__ap_idle;
  wire PEG_Bmtx_11__ap_start;
  wire PEG_Bmtx_11__ap_ready;
  wire PEG_Bmtx_11__ap_done;
  wire PEG_Bmtx_11__ap_idle;
  wire PEG_Bmtx_12__ap_start;
  wire PEG_Bmtx_12__ap_ready;
  wire PEG_Bmtx_12__ap_done;
  wire PEG_Bmtx_12__ap_idle;
  wire PEG_Bmtx_13__ap_start;
  wire PEG_Bmtx_13__ap_ready;
  wire PEG_Bmtx_13__ap_done;
  wire PEG_Bmtx_13__ap_idle;
  wire PEG_Bmtx_14__ap_start;
  wire PEG_Bmtx_14__ap_ready;
  wire PEG_Bmtx_14__ap_done;
  wire PEG_Bmtx_14__ap_idle;
  wire PEG_Bmtx_15__ap_start;
  wire PEG_Bmtx_15__ap_ready;
  wire PEG_Bmtx_15__ap_done;
  wire PEG_Bmtx_15__ap_idle;
  wire PEG_Cmtx_0__ap_start;
  wire PEG_Cmtx_0__ap_ready;
  wire PEG_Cmtx_0__ap_done;
  wire PEG_Cmtx_0__ap_idle;
  wire PEG_Cmtx_1__ap_start;
  wire PEG_Cmtx_1__ap_ready;
  wire PEG_Cmtx_1__ap_done;
  wire PEG_Cmtx_1__ap_idle;
  wire PEG_Cmtx_2__ap_start;
  wire PEG_Cmtx_2__ap_ready;
  wire PEG_Cmtx_2__ap_done;
  wire PEG_Cmtx_2__ap_idle;
  wire PEG_Cmtx_3__ap_start;
  wire PEG_Cmtx_3__ap_ready;
  wire PEG_Cmtx_3__ap_done;
  wire PEG_Cmtx_3__ap_idle;
  wire PEG_Cmtx_4__ap_start;
  wire PEG_Cmtx_4__ap_ready;
  wire PEG_Cmtx_4__ap_done;
  wire PEG_Cmtx_4__ap_idle;
  wire PEG_Cmtx_5__ap_start;
  wire PEG_Cmtx_5__ap_ready;
  wire PEG_Cmtx_5__ap_done;
  wire PEG_Cmtx_5__ap_idle;
  wire PEG_Cmtx_6__ap_start;
  wire PEG_Cmtx_6__ap_ready;
  wire PEG_Cmtx_6__ap_done;
  wire PEG_Cmtx_6__ap_idle;
  wire PEG_Cmtx_7__ap_start;
  wire PEG_Cmtx_7__ap_ready;
  wire PEG_Cmtx_7__ap_done;
  wire PEG_Cmtx_7__ap_idle;
  wire PEG_Cmtx_8__ap_start;
  wire PEG_Cmtx_8__ap_ready;
  wire PEG_Cmtx_8__ap_done;
  wire PEG_Cmtx_8__ap_idle;
  wire PEG_Cmtx_9__ap_start;
  wire PEG_Cmtx_9__ap_ready;
  wire PEG_Cmtx_9__ap_done;
  wire PEG_Cmtx_9__ap_idle;
  wire PEG_Cmtx_10__ap_start;
  wire PEG_Cmtx_10__ap_ready;
  wire PEG_Cmtx_10__ap_done;
  wire PEG_Cmtx_10__ap_idle;
  wire PEG_Cmtx_11__ap_start;
  wire PEG_Cmtx_11__ap_ready;
  wire PEG_Cmtx_11__ap_done;
  wire PEG_Cmtx_11__ap_idle;
  wire PEG_Cmtx_12__ap_start;
  wire PEG_Cmtx_12__ap_ready;
  wire PEG_Cmtx_12__ap_done;
  wire PEG_Cmtx_12__ap_idle;
  wire PEG_Cmtx_13__ap_start;
  wire PEG_Cmtx_13__ap_ready;
  wire PEG_Cmtx_13__ap_done;
  wire PEG_Cmtx_13__ap_idle;
  wire PEG_Cmtx_14__ap_start;
  wire PEG_Cmtx_14__ap_ready;
  wire PEG_Cmtx_14__ap_done;
  wire PEG_Cmtx_14__ap_idle;
  wire PEG_Cmtx_15__ap_start;
  wire PEG_Cmtx_15__ap_ready;
  wire PEG_Cmtx_15__ap_done;
  wire PEG_Cmtx_15__ap_idle;
  wire Scatter_1_2_0__ap_start;
  wire Scatter_1_2_1__ap_start;
  wire Scatter_1_2_2__ap_start;
  wire Scatter_1_2_3__ap_start;
  wire Scatter_1_2_4__ap_start;
  wire Scatter_1_2_5__ap_start;
  wire Scatter_1_2_6__ap_start;
  wire Scatter_1_2_7__ap_start;
  wire black_hole_float_v16_0__ap_start;
  wire black_hole_float_v16_1__ap_start;
  wire black_hole_float_v16_2__ap_start;
  wire black_hole_float_v16_3__ap_start;
  wire black_hole_int_0__ap_start;
  wire black_hole_int_1__ap_start;
  wire [31:0] read_A_0___NUM_A_LEN__q0;
  wire [31:0] read_A_0___P_N__q0;
  wire [63:0] read_A_0___edge_list_ch_0__q0;
  wire [63:0] edge_list_ch_0_read_addr__din;
  wire edge_list_ch_0_read_addr__full_n;
  wire edge_list_ch_0_read_addr__write;
  wire [511:0] edge_list_ch_0_read_data__dout;
  wire edge_list_ch_0_read_data__empty_n;
  wire edge_list_ch_0_read_data__read;
  wire [63:0] edge_list_ch_0_write_addr__din;
  wire edge_list_ch_0_write_addr__full_n;
  wire edge_list_ch_0_write_addr__write;
  wire [511:0] edge_list_ch_0_write_data__din;
  wire edge_list_ch_0_write_data__full_n;
  wire edge_list_ch_0_write_data__write;
  wire [7:0] edge_list_ch_0_write_resp__dout;
  wire edge_list_ch_0_write_resp__empty_n;
  wire edge_list_ch_0_write_resp__read;
  wire read_A_0__ap_start;
  wire read_A_0__ap_ready;
  wire read_A_0__ap_done;
  wire read_A_0__ap_idle;
  wire [31:0] read_A_1___NUM_A_LEN__q0;
  wire [31:0] read_A_1___P_N__q0;
  wire [63:0] read_A_1___edge_list_ch_1__q0;
  wire [63:0] edge_list_ch_1_read_addr__din;
  wire edge_list_ch_1_read_addr__full_n;
  wire edge_list_ch_1_read_addr__write;
  wire [511:0] edge_list_ch_1_read_data__dout;
  wire edge_list_ch_1_read_data__empty_n;
  wire edge_list_ch_1_read_data__read;
  wire [63:0] edge_list_ch_1_write_addr__din;
  wire edge_list_ch_1_write_addr__full_n;
  wire edge_list_ch_1_write_addr__write;
  wire [511:0] edge_list_ch_1_write_data__din;
  wire edge_list_ch_1_write_data__full_n;
  wire edge_list_ch_1_write_data__write;
  wire [7:0] edge_list_ch_1_write_resp__dout;
  wire edge_list_ch_1_write_resp__empty_n;
  wire edge_list_ch_1_write_resp__read;
  wire read_A_1__ap_start;
  wire read_A_1__ap_ready;
  wire read_A_1__ap_done;
  wire read_A_1__ap_idle;
  wire [31:0] read_A_2___NUM_A_LEN__q0;
  wire [31:0] read_A_2___P_N__q0;
  wire [63:0] read_A_2___edge_list_ch_2__q0;
  wire [63:0] edge_list_ch_2_read_addr__din;
  wire edge_list_ch_2_read_addr__full_n;
  wire edge_list_ch_2_read_addr__write;
  wire [511:0] edge_list_ch_2_read_data__dout;
  wire edge_list_ch_2_read_data__empty_n;
  wire edge_list_ch_2_read_data__read;
  wire [63:0] edge_list_ch_2_write_addr__din;
  wire edge_list_ch_2_write_addr__full_n;
  wire edge_list_ch_2_write_addr__write;
  wire [511:0] edge_list_ch_2_write_data__din;
  wire edge_list_ch_2_write_data__full_n;
  wire edge_list_ch_2_write_data__write;
  wire [7:0] edge_list_ch_2_write_resp__dout;
  wire edge_list_ch_2_write_resp__empty_n;
  wire edge_list_ch_2_write_resp__read;
  wire read_A_2__ap_start;
  wire read_A_2__ap_ready;
  wire read_A_2__ap_done;
  wire read_A_2__ap_idle;
  wire [31:0] read_A_3___NUM_A_LEN__q0;
  wire [31:0] read_A_3___P_N__q0;
  wire [63:0] read_A_3___edge_list_ch_3__q0;
  wire [63:0] edge_list_ch_3_read_addr__din;
  wire edge_list_ch_3_read_addr__full_n;
  wire edge_list_ch_3_read_addr__write;
  wire [511:0] edge_list_ch_3_read_data__dout;
  wire edge_list_ch_3_read_data__empty_n;
  wire edge_list_ch_3_read_data__read;
  wire [63:0] edge_list_ch_3_write_addr__din;
  wire edge_list_ch_3_write_addr__full_n;
  wire edge_list_ch_3_write_addr__write;
  wire [511:0] edge_list_ch_3_write_data__din;
  wire edge_list_ch_3_write_data__full_n;
  wire edge_list_ch_3_write_data__write;
  wire [7:0] edge_list_ch_3_write_resp__dout;
  wire edge_list_ch_3_write_resp__empty_n;
  wire edge_list_ch_3_write_resp__read;
  wire read_A_3__ap_start;
  wire read_A_3__ap_ready;
  wire read_A_3__ap_done;
  wire read_A_3__ap_idle;
  wire [31:0] read_A_4___NUM_A_LEN__q0;
  wire [31:0] read_A_4___P_N__q0;
  wire [63:0] read_A_4___edge_list_ch_4__q0;
  wire [63:0] edge_list_ch_4_read_addr__din;
  wire edge_list_ch_4_read_addr__full_n;
  wire edge_list_ch_4_read_addr__write;
  wire [511:0] edge_list_ch_4_read_data__dout;
  wire edge_list_ch_4_read_data__empty_n;
  wire edge_list_ch_4_read_data__read;
  wire [63:0] edge_list_ch_4_write_addr__din;
  wire edge_list_ch_4_write_addr__full_n;
  wire edge_list_ch_4_write_addr__write;
  wire [511:0] edge_list_ch_4_write_data__din;
  wire edge_list_ch_4_write_data__full_n;
  wire edge_list_ch_4_write_data__write;
  wire [7:0] edge_list_ch_4_write_resp__dout;
  wire edge_list_ch_4_write_resp__empty_n;
  wire edge_list_ch_4_write_resp__read;
  wire read_A_4__ap_start;
  wire read_A_4__ap_ready;
  wire read_A_4__ap_done;
  wire read_A_4__ap_idle;
  wire [31:0] read_A_5___NUM_A_LEN__q0;
  wire [31:0] read_A_5___P_N__q0;
  wire [63:0] read_A_5___edge_list_ch_5__q0;
  wire [63:0] edge_list_ch_5_read_addr__din;
  wire edge_list_ch_5_read_addr__full_n;
  wire edge_list_ch_5_read_addr__write;
  wire [511:0] edge_list_ch_5_read_data__dout;
  wire edge_list_ch_5_read_data__empty_n;
  wire edge_list_ch_5_read_data__read;
  wire [63:0] edge_list_ch_5_write_addr__din;
  wire edge_list_ch_5_write_addr__full_n;
  wire edge_list_ch_5_write_addr__write;
  wire [511:0] edge_list_ch_5_write_data__din;
  wire edge_list_ch_5_write_data__full_n;
  wire edge_list_ch_5_write_data__write;
  wire [7:0] edge_list_ch_5_write_resp__dout;
  wire edge_list_ch_5_write_resp__empty_n;
  wire edge_list_ch_5_write_resp__read;
  wire read_A_5__ap_start;
  wire read_A_5__ap_ready;
  wire read_A_5__ap_done;
  wire read_A_5__ap_idle;
  wire [31:0] read_A_6___NUM_A_LEN__q0;
  wire [31:0] read_A_6___P_N__q0;
  wire [63:0] read_A_6___edge_list_ch_6__q0;
  wire [63:0] edge_list_ch_6_read_addr__din;
  wire edge_list_ch_6_read_addr__full_n;
  wire edge_list_ch_6_read_addr__write;
  wire [511:0] edge_list_ch_6_read_data__dout;
  wire edge_list_ch_6_read_data__empty_n;
  wire edge_list_ch_6_read_data__read;
  wire [63:0] edge_list_ch_6_write_addr__din;
  wire edge_list_ch_6_write_addr__full_n;
  wire edge_list_ch_6_write_addr__write;
  wire [511:0] edge_list_ch_6_write_data__din;
  wire edge_list_ch_6_write_data__full_n;
  wire edge_list_ch_6_write_data__write;
  wire [7:0] edge_list_ch_6_write_resp__dout;
  wire edge_list_ch_6_write_resp__empty_n;
  wire edge_list_ch_6_write_resp__read;
  wire read_A_6__ap_start;
  wire read_A_6__ap_ready;
  wire read_A_6__ap_done;
  wire read_A_6__ap_idle;
  wire [31:0] read_A_7___NUM_A_LEN__q0;
  wire [31:0] read_A_7___P_N__q0;
  wire [63:0] read_A_7___edge_list_ch_7__q0;
  wire [63:0] edge_list_ch_7_read_addr__din;
  wire edge_list_ch_7_read_addr__full_n;
  wire edge_list_ch_7_read_addr__write;
  wire [511:0] edge_list_ch_7_read_data__dout;
  wire edge_list_ch_7_read_data__empty_n;
  wire edge_list_ch_7_read_data__read;
  wire [63:0] edge_list_ch_7_write_addr__din;
  wire edge_list_ch_7_write_addr__full_n;
  wire edge_list_ch_7_write_addr__write;
  wire [511:0] edge_list_ch_7_write_data__din;
  wire edge_list_ch_7_write_data__full_n;
  wire edge_list_ch_7_write_data__write;
  wire [7:0] edge_list_ch_7_write_resp__dout;
  wire edge_list_ch_7_write_resp__empty_n;
  wire edge_list_ch_7_write_resp__read;
  wire read_A_7__ap_start;
  wire read_A_7__ap_ready;
  wire read_A_7__ap_done;
  wire read_A_7__ap_idle;
  wire [31:0] read_B_0___K__q0;
  wire [31:0] read_B_0___P_N__q0;
  wire [63:0] read_B_0___mat_B_ch_0__q0;
  wire [63:0] mat_B_ch_0_read_addr__din;
  wire mat_B_ch_0_read_addr__full_n;
  wire mat_B_ch_0_read_addr__write;
  wire [511:0] mat_B_ch_0_read_data__dout;
  wire mat_B_ch_0_read_data__empty_n;
  wire mat_B_ch_0_read_data__read;
  wire [63:0] mat_B_ch_0_write_addr__din;
  wire mat_B_ch_0_write_addr__full_n;
  wire mat_B_ch_0_write_addr__write;
  wire [511:0] mat_B_ch_0_write_data__din;
  wire mat_B_ch_0_write_data__full_n;
  wire mat_B_ch_0_write_data__write;
  wire [7:0] mat_B_ch_0_write_resp__dout;
  wire mat_B_ch_0_write_resp__empty_n;
  wire mat_B_ch_0_write_resp__read;
  wire read_B_0__ap_start;
  wire read_B_0__ap_ready;
  wire read_B_0__ap_done;
  wire read_B_0__ap_idle;
  wire [31:0] read_B_1___K__q0;
  wire [31:0] read_B_1___P_N__q0;
  wire [63:0] read_B_1___mat_B_ch_1__q0;
  wire [63:0] mat_B_ch_1_read_addr__din;
  wire mat_B_ch_1_read_addr__full_n;
  wire mat_B_ch_1_read_addr__write;
  wire [511:0] mat_B_ch_1_read_data__dout;
  wire mat_B_ch_1_read_data__empty_n;
  wire mat_B_ch_1_read_data__read;
  wire [63:0] mat_B_ch_1_write_addr__din;
  wire mat_B_ch_1_write_addr__full_n;
  wire mat_B_ch_1_write_addr__write;
  wire [511:0] mat_B_ch_1_write_data__din;
  wire mat_B_ch_1_write_data__full_n;
  wire mat_B_ch_1_write_data__write;
  wire [7:0] mat_B_ch_1_write_resp__dout;
  wire mat_B_ch_1_write_resp__empty_n;
  wire mat_B_ch_1_write_resp__read;
  wire read_B_1__ap_start;
  wire read_B_1__ap_ready;
  wire read_B_1__ap_done;
  wire read_B_1__ap_idle;
  wire [31:0] read_B_2___K__q0;
  wire [31:0] read_B_2___P_N__q0;
  wire [63:0] read_B_2___mat_B_ch_2__q0;
  wire [63:0] mat_B_ch_2_read_addr__din;
  wire mat_B_ch_2_read_addr__full_n;
  wire mat_B_ch_2_read_addr__write;
  wire [511:0] mat_B_ch_2_read_data__dout;
  wire mat_B_ch_2_read_data__empty_n;
  wire mat_B_ch_2_read_data__read;
  wire [63:0] mat_B_ch_2_write_addr__din;
  wire mat_B_ch_2_write_addr__full_n;
  wire mat_B_ch_2_write_addr__write;
  wire [511:0] mat_B_ch_2_write_data__din;
  wire mat_B_ch_2_write_data__full_n;
  wire mat_B_ch_2_write_data__write;
  wire [7:0] mat_B_ch_2_write_resp__dout;
  wire mat_B_ch_2_write_resp__empty_n;
  wire mat_B_ch_2_write_resp__read;
  wire read_B_2__ap_start;
  wire read_B_2__ap_ready;
  wire read_B_2__ap_done;
  wire read_B_2__ap_idle;
  wire [31:0] read_B_3___K__q0;
  wire [31:0] read_B_3___P_N__q0;
  wire [63:0] read_B_3___mat_B_ch_3__q0;
  wire [63:0] mat_B_ch_3_read_addr__din;
  wire mat_B_ch_3_read_addr__full_n;
  wire mat_B_ch_3_read_addr__write;
  wire [511:0] mat_B_ch_3_read_data__dout;
  wire mat_B_ch_3_read_data__empty_n;
  wire mat_B_ch_3_read_data__read;
  wire [63:0] mat_B_ch_3_write_addr__din;
  wire mat_B_ch_3_write_addr__full_n;
  wire mat_B_ch_3_write_addr__write;
  wire [511:0] mat_B_ch_3_write_data__din;
  wire mat_B_ch_3_write_data__full_n;
  wire mat_B_ch_3_write_data__write;
  wire [7:0] mat_B_ch_3_write_resp__dout;
  wire mat_B_ch_3_write_resp__empty_n;
  wire mat_B_ch_3_write_resp__read;
  wire read_B_3__ap_start;
  wire read_B_3__ap_ready;
  wire read_B_3__ap_done;
  wire read_B_3__ap_idle;
  wire [31:0] read_C_0___M__q0;
  wire [31:0] read_C_0___P_N__q0;
  wire [63:0] read_C_0___mat_C_ch_in_0__q0;
  wire [63:0] mat_C_ch_in_0_read_addr__din;
  wire mat_C_ch_in_0_read_addr__full_n;
  wire mat_C_ch_in_0_read_addr__write;
  wire [511:0] mat_C_ch_in_0_read_data__dout;
  wire mat_C_ch_in_0_read_data__empty_n;
  wire mat_C_ch_in_0_read_data__read;
  wire [63:0] mat_C_ch_in_0_write_addr__din;
  wire mat_C_ch_in_0_write_addr__full_n;
  wire mat_C_ch_in_0_write_addr__write;
  wire [511:0] mat_C_ch_in_0_write_data__din;
  wire mat_C_ch_in_0_write_data__full_n;
  wire mat_C_ch_in_0_write_data__write;
  wire [7:0] mat_C_ch_in_0_write_resp__dout;
  wire mat_C_ch_in_0_write_resp__empty_n;
  wire mat_C_ch_in_0_write_resp__read;
  wire read_C_0__ap_start;
  wire read_C_0__ap_ready;
  wire read_C_0__ap_done;
  wire read_C_0__ap_idle;
  wire [31:0] read_C_1___M__q0;
  wire [31:0] read_C_1___P_N__q0;
  wire [63:0] read_C_1___mat_C_ch_in_1__q0;
  wire [63:0] mat_C_ch_in_1_read_addr__din;
  wire mat_C_ch_in_1_read_addr__full_n;
  wire mat_C_ch_in_1_read_addr__write;
  wire [511:0] mat_C_ch_in_1_read_data__dout;
  wire mat_C_ch_in_1_read_data__empty_n;
  wire mat_C_ch_in_1_read_data__read;
  wire [63:0] mat_C_ch_in_1_write_addr__din;
  wire mat_C_ch_in_1_write_addr__full_n;
  wire mat_C_ch_in_1_write_addr__write;
  wire [511:0] mat_C_ch_in_1_write_data__din;
  wire mat_C_ch_in_1_write_data__full_n;
  wire mat_C_ch_in_1_write_data__write;
  wire [7:0] mat_C_ch_in_1_write_resp__dout;
  wire mat_C_ch_in_1_write_resp__empty_n;
  wire mat_C_ch_in_1_write_resp__read;
  wire read_C_1__ap_start;
  wire read_C_1__ap_ready;
  wire read_C_1__ap_done;
  wire read_C_1__ap_idle;
  wire [31:0] read_C_2___M__q0;
  wire [31:0] read_C_2___P_N__q0;
  wire [63:0] read_C_2___mat_C_ch_in_2__q0;
  wire [63:0] mat_C_ch_in_2_read_addr__din;
  wire mat_C_ch_in_2_read_addr__full_n;
  wire mat_C_ch_in_2_read_addr__write;
  wire [511:0] mat_C_ch_in_2_read_data__dout;
  wire mat_C_ch_in_2_read_data__empty_n;
  wire mat_C_ch_in_2_read_data__read;
  wire [63:0] mat_C_ch_in_2_write_addr__din;
  wire mat_C_ch_in_2_write_addr__full_n;
  wire mat_C_ch_in_2_write_addr__write;
  wire [511:0] mat_C_ch_in_2_write_data__din;
  wire mat_C_ch_in_2_write_data__full_n;
  wire mat_C_ch_in_2_write_data__write;
  wire [7:0] mat_C_ch_in_2_write_resp__dout;
  wire mat_C_ch_in_2_write_resp__empty_n;
  wire mat_C_ch_in_2_write_resp__read;
  wire read_C_2__ap_start;
  wire read_C_2__ap_ready;
  wire read_C_2__ap_done;
  wire read_C_2__ap_idle;
  wire [31:0] read_C_3___M__q0;
  wire [31:0] read_C_3___P_N__q0;
  wire [63:0] read_C_3___mat_C_ch_in_3__q0;
  wire [63:0] mat_C_ch_in_3_read_addr__din;
  wire mat_C_ch_in_3_read_addr__full_n;
  wire mat_C_ch_in_3_read_addr__write;
  wire [511:0] mat_C_ch_in_3_read_data__dout;
  wire mat_C_ch_in_3_read_data__empty_n;
  wire mat_C_ch_in_3_read_data__read;
  wire [63:0] mat_C_ch_in_3_write_addr__din;
  wire mat_C_ch_in_3_write_addr__full_n;
  wire mat_C_ch_in_3_write_addr__write;
  wire [511:0] mat_C_ch_in_3_write_data__din;
  wire mat_C_ch_in_3_write_data__full_n;
  wire mat_C_ch_in_3_write_data__write;
  wire [7:0] mat_C_ch_in_3_write_resp__dout;
  wire mat_C_ch_in_3_write_resp__empty_n;
  wire mat_C_ch_in_3_write_resp__read;
  wire read_C_3__ap_start;
  wire read_C_3__ap_ready;
  wire read_C_3__ap_done;
  wire read_C_3__ap_idle;
  wire [31:0] read_C_4___M__q0;
  wire [31:0] read_C_4___P_N__q0;
  wire [63:0] read_C_4___mat_C_ch_in_4__q0;
  wire [63:0] mat_C_ch_in_4_read_addr__din;
  wire mat_C_ch_in_4_read_addr__full_n;
  wire mat_C_ch_in_4_read_addr__write;
  wire [511:0] mat_C_ch_in_4_read_data__dout;
  wire mat_C_ch_in_4_read_data__empty_n;
  wire mat_C_ch_in_4_read_data__read;
  wire [63:0] mat_C_ch_in_4_write_addr__din;
  wire mat_C_ch_in_4_write_addr__full_n;
  wire mat_C_ch_in_4_write_addr__write;
  wire [511:0] mat_C_ch_in_4_write_data__din;
  wire mat_C_ch_in_4_write_data__full_n;
  wire mat_C_ch_in_4_write_data__write;
  wire [7:0] mat_C_ch_in_4_write_resp__dout;
  wire mat_C_ch_in_4_write_resp__empty_n;
  wire mat_C_ch_in_4_write_resp__read;
  wire read_C_4__ap_start;
  wire read_C_4__ap_ready;
  wire read_C_4__ap_done;
  wire read_C_4__ap_idle;
  wire [31:0] read_C_5___M__q0;
  wire [31:0] read_C_5___P_N__q0;
  wire [63:0] read_C_5___mat_C_ch_in_5__q0;
  wire [63:0] mat_C_ch_in_5_read_addr__din;
  wire mat_C_ch_in_5_read_addr__full_n;
  wire mat_C_ch_in_5_read_addr__write;
  wire [511:0] mat_C_ch_in_5_read_data__dout;
  wire mat_C_ch_in_5_read_data__empty_n;
  wire mat_C_ch_in_5_read_data__read;
  wire [63:0] mat_C_ch_in_5_write_addr__din;
  wire mat_C_ch_in_5_write_addr__full_n;
  wire mat_C_ch_in_5_write_addr__write;
  wire [511:0] mat_C_ch_in_5_write_data__din;
  wire mat_C_ch_in_5_write_data__full_n;
  wire mat_C_ch_in_5_write_data__write;
  wire [7:0] mat_C_ch_in_5_write_resp__dout;
  wire mat_C_ch_in_5_write_resp__empty_n;
  wire mat_C_ch_in_5_write_resp__read;
  wire read_C_5__ap_start;
  wire read_C_5__ap_ready;
  wire read_C_5__ap_done;
  wire read_C_5__ap_idle;
  wire [31:0] read_C_6___M__q0;
  wire [31:0] read_C_6___P_N__q0;
  wire [63:0] read_C_6___mat_C_ch_in_6__q0;
  wire [63:0] mat_C_ch_in_6_read_addr__din;
  wire mat_C_ch_in_6_read_addr__full_n;
  wire mat_C_ch_in_6_read_addr__write;
  wire [511:0] mat_C_ch_in_6_read_data__dout;
  wire mat_C_ch_in_6_read_data__empty_n;
  wire mat_C_ch_in_6_read_data__read;
  wire [63:0] mat_C_ch_in_6_write_addr__din;
  wire mat_C_ch_in_6_write_addr__full_n;
  wire mat_C_ch_in_6_write_addr__write;
  wire [511:0] mat_C_ch_in_6_write_data__din;
  wire mat_C_ch_in_6_write_data__full_n;
  wire mat_C_ch_in_6_write_data__write;
  wire [7:0] mat_C_ch_in_6_write_resp__dout;
  wire mat_C_ch_in_6_write_resp__empty_n;
  wire mat_C_ch_in_6_write_resp__read;
  wire read_C_6__ap_start;
  wire read_C_6__ap_ready;
  wire read_C_6__ap_done;
  wire read_C_6__ap_idle;
  wire [31:0] read_C_7___M__q0;
  wire [31:0] read_C_7___P_N__q0;
  wire [63:0] read_C_7___mat_C_ch_in_7__q0;
  wire [63:0] mat_C_ch_in_7_read_addr__din;
  wire mat_C_ch_in_7_read_addr__full_n;
  wire mat_C_ch_in_7_read_addr__write;
  wire [511:0] mat_C_ch_in_7_read_data__dout;
  wire mat_C_ch_in_7_read_data__empty_n;
  wire mat_C_ch_in_7_read_data__read;
  wire [63:0] mat_C_ch_in_7_write_addr__din;
  wire mat_C_ch_in_7_write_addr__full_n;
  wire mat_C_ch_in_7_write_addr__write;
  wire [511:0] mat_C_ch_in_7_write_data__din;
  wire mat_C_ch_in_7_write_data__full_n;
  wire mat_C_ch_in_7_write_data__write;
  wire [7:0] mat_C_ch_in_7_write_resp__dout;
  wire mat_C_ch_in_7_write_resp__empty_n;
  wire mat_C_ch_in_7_write_resp__read;
  wire read_C_7__ap_start;
  wire read_C_7__ap_ready;
  wire read_C_7__ap_done;
  wire read_C_7__ap_idle;
  wire [31:0] read_edge_list_ptr_0___K__q0;
  wire [31:0] read_edge_list_ptr_0___M__q0;
  wire [31:0] read_edge_list_ptr_0___NUM_ITE__q0;
  wire [31:0] read_edge_list_ptr_0___P_N__q0;
  wire [63:0] read_edge_list_ptr_0___edge_list_ptr__q0;
  wire [63:0] edge_list_ptr_read_addr__din;
  wire edge_list_ptr_read_addr__full_n;
  wire edge_list_ptr_read_addr__write;
  wire [31:0] edge_list_ptr_read_data__dout;
  wire edge_list_ptr_read_data__empty_n;
  wire edge_list_ptr_read_data__read;
  wire [63:0] edge_list_ptr_write_addr__din;
  wire edge_list_ptr_write_addr__full_n;
  wire edge_list_ptr_write_addr__write;
  wire [31:0] edge_list_ptr_write_data__din;
  wire edge_list_ptr_write_data__full_n;
  wire edge_list_ptr_write_data__write;
  wire [7:0] edge_list_ptr_write_resp__dout;
  wire edge_list_ptr_write_resp__empty_n;
  wire edge_list_ptr_write_resp__read;
  wire read_edge_list_ptr_0__ap_start;
  wire read_edge_list_ptr_0__ap_ready;
  wire read_edge_list_ptr_0__ap_done;
  wire read_edge_list_ptr_0__ap_idle;
  wire [63:0] write_C_0___mat_C_ch_0__q0;
  wire [63:0] mat_C_ch_0_read_addr__din;
  wire mat_C_ch_0_read_addr__full_n;
  wire mat_C_ch_0_read_addr__write;
  wire [511:0] mat_C_ch_0_read_data__dout;
  wire mat_C_ch_0_read_data__empty_n;
  wire mat_C_ch_0_read_data__read;
  wire [63:0] mat_C_ch_0_write_addr__din;
  wire mat_C_ch_0_write_addr__full_n;
  wire mat_C_ch_0_write_addr__write;
  wire [511:0] mat_C_ch_0_write_data__din;
  wire mat_C_ch_0_write_data__full_n;
  wire mat_C_ch_0_write_data__write;
  wire [7:0] mat_C_ch_0_write_resp__dout;
  wire mat_C_ch_0_write_resp__empty_n;
  wire mat_C_ch_0_write_resp__read;
  wire write_C_0__ap_start;
  wire write_C_0__ap_ready;
  wire write_C_0__ap_done;
  wire write_C_0__ap_idle;
  wire [63:0] write_C_1___mat_C_ch_1__q0;
  wire [63:0] mat_C_ch_1_read_addr__din;
  wire mat_C_ch_1_read_addr__full_n;
  wire mat_C_ch_1_read_addr__write;
  wire [511:0] mat_C_ch_1_read_data__dout;
  wire mat_C_ch_1_read_data__empty_n;
  wire mat_C_ch_1_read_data__read;
  wire [63:0] mat_C_ch_1_write_addr__din;
  wire mat_C_ch_1_write_addr__full_n;
  wire mat_C_ch_1_write_addr__write;
  wire [511:0] mat_C_ch_1_write_data__din;
  wire mat_C_ch_1_write_data__full_n;
  wire mat_C_ch_1_write_data__write;
  wire [7:0] mat_C_ch_1_write_resp__dout;
  wire mat_C_ch_1_write_resp__empty_n;
  wire mat_C_ch_1_write_resp__read;
  wire write_C_1__ap_start;
  wire write_C_1__ap_ready;
  wire write_C_1__ap_done;
  wire write_C_1__ap_idle;
  wire [63:0] write_C_2___mat_C_ch_2__q0;
  wire [63:0] mat_C_ch_2_read_addr__din;
  wire mat_C_ch_2_read_addr__full_n;
  wire mat_C_ch_2_read_addr__write;
  wire [511:0] mat_C_ch_2_read_data__dout;
  wire mat_C_ch_2_read_data__empty_n;
  wire mat_C_ch_2_read_data__read;
  wire [63:0] mat_C_ch_2_write_addr__din;
  wire mat_C_ch_2_write_addr__full_n;
  wire mat_C_ch_2_write_addr__write;
  wire [511:0] mat_C_ch_2_write_data__din;
  wire mat_C_ch_2_write_data__full_n;
  wire mat_C_ch_2_write_data__write;
  wire [7:0] mat_C_ch_2_write_resp__dout;
  wire mat_C_ch_2_write_resp__empty_n;
  wire mat_C_ch_2_write_resp__read;
  wire write_C_2__ap_start;
  wire write_C_2__ap_ready;
  wire write_C_2__ap_done;
  wire write_C_2__ap_idle;
  wire [63:0] write_C_3___mat_C_ch_3__q0;
  wire [63:0] mat_C_ch_3_read_addr__din;
  wire mat_C_ch_3_read_addr__full_n;
  wire mat_C_ch_3_read_addr__write;
  wire [511:0] mat_C_ch_3_read_data__dout;
  wire mat_C_ch_3_read_data__empty_n;
  wire mat_C_ch_3_read_data__read;
  wire [63:0] mat_C_ch_3_write_addr__din;
  wire mat_C_ch_3_write_addr__full_n;
  wire mat_C_ch_3_write_addr__write;
  wire [511:0] mat_C_ch_3_write_data__din;
  wire mat_C_ch_3_write_data__full_n;
  wire mat_C_ch_3_write_data__write;
  wire [7:0] mat_C_ch_3_write_resp__dout;
  wire mat_C_ch_3_write_resp__empty_n;
  wire mat_C_ch_3_write_resp__read;
  wire write_C_3__ap_start;
  wire write_C_3__ap_ready;
  wire write_C_3__ap_done;
  wire write_C_3__ap_idle;
  wire [63:0] write_C_4___mat_C_ch_4__q0;
  wire [63:0] mat_C_ch_4_read_addr__din;
  wire mat_C_ch_4_read_addr__full_n;
  wire mat_C_ch_4_read_addr__write;
  wire [511:0] mat_C_ch_4_read_data__dout;
  wire mat_C_ch_4_read_data__empty_n;
  wire mat_C_ch_4_read_data__read;
  wire [63:0] mat_C_ch_4_write_addr__din;
  wire mat_C_ch_4_write_addr__full_n;
  wire mat_C_ch_4_write_addr__write;
  wire [511:0] mat_C_ch_4_write_data__din;
  wire mat_C_ch_4_write_data__full_n;
  wire mat_C_ch_4_write_data__write;
  wire [7:0] mat_C_ch_4_write_resp__dout;
  wire mat_C_ch_4_write_resp__empty_n;
  wire mat_C_ch_4_write_resp__read;
  wire write_C_4__ap_start;
  wire write_C_4__ap_ready;
  wire write_C_4__ap_done;
  wire write_C_4__ap_idle;
  wire [63:0] write_C_5___mat_C_ch_5__q0;
  wire [63:0] mat_C_ch_5_read_addr__din;
  wire mat_C_ch_5_read_addr__full_n;
  wire mat_C_ch_5_read_addr__write;
  wire [511:0] mat_C_ch_5_read_data__dout;
  wire mat_C_ch_5_read_data__empty_n;
  wire mat_C_ch_5_read_data__read;
  wire [63:0] mat_C_ch_5_write_addr__din;
  wire mat_C_ch_5_write_addr__full_n;
  wire mat_C_ch_5_write_addr__write;
  wire [511:0] mat_C_ch_5_write_data__din;
  wire mat_C_ch_5_write_data__full_n;
  wire mat_C_ch_5_write_data__write;
  wire [7:0] mat_C_ch_5_write_resp__dout;
  wire mat_C_ch_5_write_resp__empty_n;
  wire mat_C_ch_5_write_resp__read;
  wire write_C_5__ap_start;
  wire write_C_5__ap_ready;
  wire write_C_5__ap_done;
  wire write_C_5__ap_idle;
  wire [63:0] write_C_6___mat_C_ch_6__q0;
  wire [63:0] mat_C_ch_6_read_addr__din;
  wire mat_C_ch_6_read_addr__full_n;
  wire mat_C_ch_6_read_addr__write;
  wire [511:0] mat_C_ch_6_read_data__dout;
  wire mat_C_ch_6_read_data__empty_n;
  wire mat_C_ch_6_read_data__read;
  wire [63:0] mat_C_ch_6_write_addr__din;
  wire mat_C_ch_6_write_addr__full_n;
  wire mat_C_ch_6_write_addr__write;
  wire [511:0] mat_C_ch_6_write_data__din;
  wire mat_C_ch_6_write_data__full_n;
  wire mat_C_ch_6_write_data__write;
  wire [7:0] mat_C_ch_6_write_resp__dout;
  wire mat_C_ch_6_write_resp__empty_n;
  wire mat_C_ch_6_write_resp__read;
  wire write_C_6__ap_start;
  wire write_C_6__ap_ready;
  wire write_C_6__ap_done;
  wire write_C_6__ap_idle;
  wire [63:0] write_C_7___mat_C_ch_7__q0;
  wire [63:0] mat_C_ch_7_read_addr__din;
  wire mat_C_ch_7_read_addr__full_n;
  wire mat_C_ch_7_read_addr__write;
  wire [511:0] mat_C_ch_7_read_data__dout;
  wire mat_C_ch_7_read_data__empty_n;
  wire mat_C_ch_7_read_data__read;
  wire [63:0] mat_C_ch_7_write_addr__din;
  wire mat_C_ch_7_write_addr__full_n;
  wire mat_C_ch_7_write_addr__write;
  wire [511:0] mat_C_ch_7_write_data__din;
  wire mat_C_ch_7_write_data__full_n;
  wire mat_C_ch_7_write_data__write;
  wire [7:0] mat_C_ch_7_write_resp__dout;
  wire mat_C_ch_7_write_resp__empty_n;
  wire mat_C_ch_7_write_resp__read;
  wire write_C_7__ap_start;
  wire write_C_7__ap_ready;
  wire write_C_7__ap_done;
  wire write_C_7__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;

  Sextans_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .edge_list_ptr(edge_list_ptr),
    .edge_list_ch_0(edge_list_ch_0),
    .edge_list_ch_1(edge_list_ch_1),
    .edge_list_ch_2(edge_list_ch_2),
    .edge_list_ch_3(edge_list_ch_3),
    .edge_list_ch_4(edge_list_ch_4),
    .edge_list_ch_5(edge_list_ch_5),
    .edge_list_ch_6(edge_list_ch_6),
    .edge_list_ch_7(edge_list_ch_7),
    .mat_B_ch_0(mat_B_ch_0),
    .mat_B_ch_1(mat_B_ch_1),
    .mat_B_ch_2(mat_B_ch_2),
    .mat_B_ch_3(mat_B_ch_3),
    .mat_C_ch_in_0(mat_C_ch_in_0),
    .mat_C_ch_in_1(mat_C_ch_in_1),
    .mat_C_ch_in_2(mat_C_ch_in_2),
    .mat_C_ch_in_3(mat_C_ch_in_3),
    .mat_C_ch_in_4(mat_C_ch_in_4),
    .mat_C_ch_in_5(mat_C_ch_in_5),
    .mat_C_ch_in_6(mat_C_ch_in_6),
    .mat_C_ch_in_7(mat_C_ch_in_7),
    .mat_C_ch_0(mat_C_ch_0),
    .mat_C_ch_1(mat_C_ch_1),
    .mat_C_ch_2(mat_C_ch_2),
    .mat_C_ch_3(mat_C_ch_3),
    .mat_C_ch_4(mat_C_ch_4),
    .mat_C_ch_5(mat_C_ch_5),
    .mat_C_ch_6(mat_C_ch_6),
    .mat_C_ch_7(mat_C_ch_7),
    .NUM_ITE(NUM_ITE),
    .NUM_A_LEN(NUM_A_LEN),
    .M(M),
    .K(K),
    .P_N(P_N),
    .alpha_u(alpha_u),
    .beta_u(beta_u),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_0__dout),
    .if_empty_n(PE_inst_Sextans_0__empty_n),
    .if_read(PE_inst_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_0__din),
    .if_full_n(PE_inst_Sextans_0__full_n),
    .if_write(PE_inst_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_10__dout),
    .if_empty_n(PE_inst_Sextans_10__empty_n),
    .if_read(PE_inst_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_10__din),
    .if_full_n(PE_inst_Sextans_10__full_n),
    .if_write(PE_inst_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_11__dout),
    .if_empty_n(PE_inst_Sextans_11__empty_n),
    .if_read(PE_inst_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_11__din),
    .if_full_n(PE_inst_Sextans_11__full_n),
    .if_write(PE_inst_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_12__dout),
    .if_empty_n(PE_inst_Sextans_12__empty_n),
    .if_read(PE_inst_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_12__din),
    .if_full_n(PE_inst_Sextans_12__full_n),
    .if_write(PE_inst_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_13__dout),
    .if_empty_n(PE_inst_Sextans_13__empty_n),
    .if_read(PE_inst_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_13__din),
    .if_full_n(PE_inst_Sextans_13__full_n),
    .if_write(PE_inst_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_14__dout),
    .if_empty_n(PE_inst_Sextans_14__empty_n),
    .if_read(PE_inst_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_14__din),
    .if_full_n(PE_inst_Sextans_14__full_n),
    .if_write(PE_inst_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_15__dout),
    .if_empty_n(PE_inst_Sextans_15__empty_n),
    .if_read(PE_inst_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_15__din),
    .if_full_n(PE_inst_Sextans_15__full_n),
    .if_write(PE_inst_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_16__dout),
    .if_empty_n(PE_inst_Sextans_16__empty_n),
    .if_read(PE_inst_Sextans_16__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_16__din),
    .if_full_n(PE_inst_Sextans_16__full_n),
    .if_write(PE_inst_Sextans_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_1__dout),
    .if_empty_n(PE_inst_Sextans_1__empty_n),
    .if_read(PE_inst_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_1__din),
    .if_full_n(PE_inst_Sextans_1__full_n),
    .if_write(PE_inst_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_2__dout),
    .if_empty_n(PE_inst_Sextans_2__empty_n),
    .if_read(PE_inst_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_2__din),
    .if_full_n(PE_inst_Sextans_2__full_n),
    .if_write(PE_inst_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_3__dout),
    .if_empty_n(PE_inst_Sextans_3__empty_n),
    .if_read(PE_inst_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_3__din),
    .if_full_n(PE_inst_Sextans_3__full_n),
    .if_write(PE_inst_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_4__dout),
    .if_empty_n(PE_inst_Sextans_4__empty_n),
    .if_read(PE_inst_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_4__din),
    .if_full_n(PE_inst_Sextans_4__full_n),
    .if_write(PE_inst_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_5__dout),
    .if_empty_n(PE_inst_Sextans_5__empty_n),
    .if_read(PE_inst_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_5__din),
    .if_full_n(PE_inst_Sextans_5__full_n),
    .if_write(PE_inst_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_6__dout),
    .if_empty_n(PE_inst_Sextans_6__empty_n),
    .if_read(PE_inst_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_6__din),
    .if_full_n(PE_inst_Sextans_6__full_n),
    .if_write(PE_inst_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_7__dout),
    .if_empty_n(PE_inst_Sextans_7__empty_n),
    .if_read(PE_inst_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_7__din),
    .if_full_n(PE_inst_Sextans_7__full_n),
    .if_write(PE_inst_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_8__dout),
    .if_empty_n(PE_inst_Sextans_8__empty_n),
    .if_read(PE_inst_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_8__din),
    .if_full_n(PE_inst_Sextans_8__full_n),
    .if_write(PE_inst_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_Sextans_9__dout),
    .if_empty_n(PE_inst_Sextans_9__empty_n),
    .if_read(PE_inst_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_Sextans_9__din),
    .if_full_n(PE_inst_Sextans_9__full_n),
    .if_write(PE_inst_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_0__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_0__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_0__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_0__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_10__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_10__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_10__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_10__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_11__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_11__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_11__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_11__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_12__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_12__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_12__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_12__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_13__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_13__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_13__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_13__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_14__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_14__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_14__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_14__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_15__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_15__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_15__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_15__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_1__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_1__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_1__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_1__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_2__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_2__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_2__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_2__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_3__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_3__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_3__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_3__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_4__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_4__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_4__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_4__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_5__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_5__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_5__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_5__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_6__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_6__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_6__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_6__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_7__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_7__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_7__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_7__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_8__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_8__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_8__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_8__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  PE_inst_to_Cmtx_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(PE_inst_to_Cmtx_Sextans_9__dout),
    .if_empty_n(PE_inst_to_Cmtx_Sextans_9__empty_n),
    .if_read(PE_inst_to_Cmtx_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(PE_inst_to_Cmtx_Sextans_9__din),
    .if_full_n(PE_inst_to_Cmtx_Sextans_9__full_n),
    .if_write(PE_inst_to_Cmtx_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_0__dout),
    .if_empty_n(fifo_A_Sextans_0__empty_n),
    .if_read(fifo_A_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_0__din),
    .if_full_n(fifo_A_Sextans_0__full_n),
    .if_write(fifo_A_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_1__dout),
    .if_empty_n(fifo_A_Sextans_1__empty_n),
    .if_read(fifo_A_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_1__din),
    .if_full_n(fifo_A_Sextans_1__full_n),
    .if_write(fifo_A_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_2__dout),
    .if_empty_n(fifo_A_Sextans_2__empty_n),
    .if_read(fifo_A_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_2__din),
    .if_full_n(fifo_A_Sextans_2__full_n),
    .if_write(fifo_A_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_3__dout),
    .if_empty_n(fifo_A_Sextans_3__empty_n),
    .if_read(fifo_A_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_3__din),
    .if_full_n(fifo_A_Sextans_3__full_n),
    .if_write(fifo_A_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_4__dout),
    .if_empty_n(fifo_A_Sextans_4__empty_n),
    .if_read(fifo_A_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_4__din),
    .if_full_n(fifo_A_Sextans_4__full_n),
    .if_write(fifo_A_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_5__dout),
    .if_empty_n(fifo_A_Sextans_5__empty_n),
    .if_read(fifo_A_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_5__din),
    .if_full_n(fifo_A_Sextans_5__full_n),
    .if_write(fifo_A_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_6__dout),
    .if_empty_n(fifo_A_Sextans_6__empty_n),
    .if_read(fifo_A_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_6__din),
    .if_full_n(fifo_A_Sextans_6__full_n),
    .if_write(fifo_A_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_Sextans_7__dout),
    .if_empty_n(fifo_A_Sextans_7__empty_n),
    .if_read(fifo_A_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_Sextans_7__din),
    .if_full_n(fifo_A_Sextans_7__full_n),
    .if_write(fifo_A_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_0__dout),
    .if_empty_n(fifo_A_pe_Sextans_0__empty_n),
    .if_read(fifo_A_pe_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_0__din),
    .if_full_n(fifo_A_pe_Sextans_0__full_n),
    .if_write(fifo_A_pe_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_10__dout),
    .if_empty_n(fifo_A_pe_Sextans_10__empty_n),
    .if_read(fifo_A_pe_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_10__din),
    .if_full_n(fifo_A_pe_Sextans_10__full_n),
    .if_write(fifo_A_pe_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_11__dout),
    .if_empty_n(fifo_A_pe_Sextans_11__empty_n),
    .if_read(fifo_A_pe_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_11__din),
    .if_full_n(fifo_A_pe_Sextans_11__full_n),
    .if_write(fifo_A_pe_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_12__dout),
    .if_empty_n(fifo_A_pe_Sextans_12__empty_n),
    .if_read(fifo_A_pe_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_12__din),
    .if_full_n(fifo_A_pe_Sextans_12__full_n),
    .if_write(fifo_A_pe_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_13__dout),
    .if_empty_n(fifo_A_pe_Sextans_13__empty_n),
    .if_read(fifo_A_pe_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_13__din),
    .if_full_n(fifo_A_pe_Sextans_13__full_n),
    .if_write(fifo_A_pe_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_14__dout),
    .if_empty_n(fifo_A_pe_Sextans_14__empty_n),
    .if_read(fifo_A_pe_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_14__din),
    .if_full_n(fifo_A_pe_Sextans_14__full_n),
    .if_write(fifo_A_pe_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_15__dout),
    .if_empty_n(fifo_A_pe_Sextans_15__empty_n),
    .if_read(fifo_A_pe_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_15__din),
    .if_full_n(fifo_A_pe_Sextans_15__full_n),
    .if_write(fifo_A_pe_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_1__dout),
    .if_empty_n(fifo_A_pe_Sextans_1__empty_n),
    .if_read(fifo_A_pe_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_1__din),
    .if_full_n(fifo_A_pe_Sextans_1__full_n),
    .if_write(fifo_A_pe_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_2__dout),
    .if_empty_n(fifo_A_pe_Sextans_2__empty_n),
    .if_read(fifo_A_pe_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_2__din),
    .if_full_n(fifo_A_pe_Sextans_2__full_n),
    .if_write(fifo_A_pe_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_3__dout),
    .if_empty_n(fifo_A_pe_Sextans_3__empty_n),
    .if_read(fifo_A_pe_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_3__din),
    .if_full_n(fifo_A_pe_Sextans_3__full_n),
    .if_write(fifo_A_pe_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_4__dout),
    .if_empty_n(fifo_A_pe_Sextans_4__empty_n),
    .if_read(fifo_A_pe_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_4__din),
    .if_full_n(fifo_A_pe_Sextans_4__full_n),
    .if_write(fifo_A_pe_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_5__dout),
    .if_empty_n(fifo_A_pe_Sextans_5__empty_n),
    .if_read(fifo_A_pe_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_5__din),
    .if_full_n(fifo_A_pe_Sextans_5__full_n),
    .if_write(fifo_A_pe_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_6__dout),
    .if_empty_n(fifo_A_pe_Sextans_6__empty_n),
    .if_read(fifo_A_pe_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_6__din),
    .if_full_n(fifo_A_pe_Sextans_6__full_n),
    .if_write(fifo_A_pe_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_7__dout),
    .if_empty_n(fifo_A_pe_Sextans_7__empty_n),
    .if_read(fifo_A_pe_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_7__din),
    .if_full_n(fifo_A_pe_Sextans_7__full_n),
    .if_write(fifo_A_pe_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_8__dout),
    .if_empty_n(fifo_A_pe_Sextans_8__empty_n),
    .if_read(fifo_A_pe_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_8__din),
    .if_full_n(fifo_A_pe_Sextans_8__full_n),
    .if_write(fifo_A_pe_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_pe_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_pe_Sextans_9__dout),
    .if_empty_n(fifo_A_pe_Sextans_9__empty_n),
    .if_read(fifo_A_pe_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_pe_Sextans_9__din),
    .if_full_n(fifo_A_pe_Sextans_9__full_n),
    .if_write(fifo_A_pe_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_0__dout),
    .if_empty_n(fifo_B_pe_Sextans_0__empty_n),
    .if_read(fifo_B_pe_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_0__din),
    .if_full_n(fifo_B_pe_Sextans_0__full_n),
    .if_write(fifo_B_pe_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_10__dout),
    .if_empty_n(fifo_B_pe_Sextans_10__empty_n),
    .if_read(fifo_B_pe_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_10__din),
    .if_full_n(fifo_B_pe_Sextans_10__full_n),
    .if_write(fifo_B_pe_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_11__dout),
    .if_empty_n(fifo_B_pe_Sextans_11__empty_n),
    .if_read(fifo_B_pe_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_11__din),
    .if_full_n(fifo_B_pe_Sextans_11__full_n),
    .if_write(fifo_B_pe_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_12__dout),
    .if_empty_n(fifo_B_pe_Sextans_12__empty_n),
    .if_read(fifo_B_pe_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_12__din),
    .if_full_n(fifo_B_pe_Sextans_12__full_n),
    .if_write(fifo_B_pe_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_13__dout),
    .if_empty_n(fifo_B_pe_Sextans_13__empty_n),
    .if_read(fifo_B_pe_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_13__din),
    .if_full_n(fifo_B_pe_Sextans_13__full_n),
    .if_write(fifo_B_pe_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_14__dout),
    .if_empty_n(fifo_B_pe_Sextans_14__empty_n),
    .if_read(fifo_B_pe_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_14__din),
    .if_full_n(fifo_B_pe_Sextans_14__full_n),
    .if_write(fifo_B_pe_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_15__dout),
    .if_empty_n(fifo_B_pe_Sextans_15__empty_n),
    .if_read(fifo_B_pe_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_15__din),
    .if_full_n(fifo_B_pe_Sextans_15__full_n),
    .if_write(fifo_B_pe_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_16__dout),
    .if_empty_n(fifo_B_pe_Sextans_16__empty_n),
    .if_read(fifo_B_pe_Sextans_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_16__din),
    .if_full_n(fifo_B_pe_Sextans_16__full_n),
    .if_write(fifo_B_pe_Sextans_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_17__dout),
    .if_empty_n(fifo_B_pe_Sextans_17__empty_n),
    .if_read(fifo_B_pe_Sextans_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_17__din),
    .if_full_n(fifo_B_pe_Sextans_17__full_n),
    .if_write(fifo_B_pe_Sextans_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_18
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_18__dout),
    .if_empty_n(fifo_B_pe_Sextans_18__empty_n),
    .if_read(fifo_B_pe_Sextans_18__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_18__din),
    .if_full_n(fifo_B_pe_Sextans_18__full_n),
    .if_write(fifo_B_pe_Sextans_18__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_19
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_19__dout),
    .if_empty_n(fifo_B_pe_Sextans_19__empty_n),
    .if_read(fifo_B_pe_Sextans_19__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_19__din),
    .if_full_n(fifo_B_pe_Sextans_19__full_n),
    .if_write(fifo_B_pe_Sextans_19__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_1__dout),
    .if_empty_n(fifo_B_pe_Sextans_1__empty_n),
    .if_read(fifo_B_pe_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_1__din),
    .if_full_n(fifo_B_pe_Sextans_1__full_n),
    .if_write(fifo_B_pe_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_20
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_20__dout),
    .if_empty_n(fifo_B_pe_Sextans_20__empty_n),
    .if_read(fifo_B_pe_Sextans_20__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_20__din),
    .if_full_n(fifo_B_pe_Sextans_20__full_n),
    .if_write(fifo_B_pe_Sextans_20__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_21
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_21__dout),
    .if_empty_n(fifo_B_pe_Sextans_21__empty_n),
    .if_read(fifo_B_pe_Sextans_21__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_21__din),
    .if_full_n(fifo_B_pe_Sextans_21__full_n),
    .if_write(fifo_B_pe_Sextans_21__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_22
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_22__dout),
    .if_empty_n(fifo_B_pe_Sextans_22__empty_n),
    .if_read(fifo_B_pe_Sextans_22__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_22__din),
    .if_full_n(fifo_B_pe_Sextans_22__full_n),
    .if_write(fifo_B_pe_Sextans_22__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_23
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_23__dout),
    .if_empty_n(fifo_B_pe_Sextans_23__empty_n),
    .if_read(fifo_B_pe_Sextans_23__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_23__din),
    .if_full_n(fifo_B_pe_Sextans_23__full_n),
    .if_write(fifo_B_pe_Sextans_23__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_24
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_24__dout),
    .if_empty_n(fifo_B_pe_Sextans_24__empty_n),
    .if_read(fifo_B_pe_Sextans_24__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_24__din),
    .if_full_n(fifo_B_pe_Sextans_24__full_n),
    .if_write(fifo_B_pe_Sextans_24__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_25
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_25__dout),
    .if_empty_n(fifo_B_pe_Sextans_25__empty_n),
    .if_read(fifo_B_pe_Sextans_25__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_25__din),
    .if_full_n(fifo_B_pe_Sextans_25__full_n),
    .if_write(fifo_B_pe_Sextans_25__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_26
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_26__dout),
    .if_empty_n(fifo_B_pe_Sextans_26__empty_n),
    .if_read(fifo_B_pe_Sextans_26__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_26__din),
    .if_full_n(fifo_B_pe_Sextans_26__full_n),
    .if_write(fifo_B_pe_Sextans_26__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_27
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_27__dout),
    .if_empty_n(fifo_B_pe_Sextans_27__empty_n),
    .if_read(fifo_B_pe_Sextans_27__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_27__din),
    .if_full_n(fifo_B_pe_Sextans_27__full_n),
    .if_write(fifo_B_pe_Sextans_27__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_28
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_28__dout),
    .if_empty_n(fifo_B_pe_Sextans_28__empty_n),
    .if_read(fifo_B_pe_Sextans_28__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_28__din),
    .if_full_n(fifo_B_pe_Sextans_28__full_n),
    .if_write(fifo_B_pe_Sextans_28__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_29
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_29__dout),
    .if_empty_n(fifo_B_pe_Sextans_29__empty_n),
    .if_read(fifo_B_pe_Sextans_29__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_29__din),
    .if_full_n(fifo_B_pe_Sextans_29__full_n),
    .if_write(fifo_B_pe_Sextans_29__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_2__dout),
    .if_empty_n(fifo_B_pe_Sextans_2__empty_n),
    .if_read(fifo_B_pe_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_2__din),
    .if_full_n(fifo_B_pe_Sextans_2__full_n),
    .if_write(fifo_B_pe_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_30
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_30__dout),
    .if_empty_n(fifo_B_pe_Sextans_30__empty_n),
    .if_read(fifo_B_pe_Sextans_30__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_30__din),
    .if_full_n(fifo_B_pe_Sextans_30__full_n),
    .if_write(fifo_B_pe_Sextans_30__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_31
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_31__dout),
    .if_empty_n(fifo_B_pe_Sextans_31__empty_n),
    .if_read(fifo_B_pe_Sextans_31__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_31__din),
    .if_full_n(fifo_B_pe_Sextans_31__full_n),
    .if_write(fifo_B_pe_Sextans_31__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_32
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_32__dout),
    .if_empty_n(fifo_B_pe_Sextans_32__empty_n),
    .if_read(fifo_B_pe_Sextans_32__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_32__din),
    .if_full_n(fifo_B_pe_Sextans_32__full_n),
    .if_write(fifo_B_pe_Sextans_32__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_33
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_33__dout),
    .if_empty_n(fifo_B_pe_Sextans_33__empty_n),
    .if_read(fifo_B_pe_Sextans_33__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_33__din),
    .if_full_n(fifo_B_pe_Sextans_33__full_n),
    .if_write(fifo_B_pe_Sextans_33__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_34
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_34__dout),
    .if_empty_n(fifo_B_pe_Sextans_34__empty_n),
    .if_read(fifo_B_pe_Sextans_34__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_34__din),
    .if_full_n(fifo_B_pe_Sextans_34__full_n),
    .if_write(fifo_B_pe_Sextans_34__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_35
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_35__dout),
    .if_empty_n(fifo_B_pe_Sextans_35__empty_n),
    .if_read(fifo_B_pe_Sextans_35__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_35__din),
    .if_full_n(fifo_B_pe_Sextans_35__full_n),
    .if_write(fifo_B_pe_Sextans_35__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_36
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_36__dout),
    .if_empty_n(fifo_B_pe_Sextans_36__empty_n),
    .if_read(fifo_B_pe_Sextans_36__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_36__din),
    .if_full_n(fifo_B_pe_Sextans_36__full_n),
    .if_write(fifo_B_pe_Sextans_36__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_37
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_37__dout),
    .if_empty_n(fifo_B_pe_Sextans_37__empty_n),
    .if_read(fifo_B_pe_Sextans_37__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_37__din),
    .if_full_n(fifo_B_pe_Sextans_37__full_n),
    .if_write(fifo_B_pe_Sextans_37__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_38
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_38__dout),
    .if_empty_n(fifo_B_pe_Sextans_38__empty_n),
    .if_read(fifo_B_pe_Sextans_38__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_38__din),
    .if_full_n(fifo_B_pe_Sextans_38__full_n),
    .if_write(fifo_B_pe_Sextans_38__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_39
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_39__dout),
    .if_empty_n(fifo_B_pe_Sextans_39__empty_n),
    .if_read(fifo_B_pe_Sextans_39__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_39__din),
    .if_full_n(fifo_B_pe_Sextans_39__full_n),
    .if_write(fifo_B_pe_Sextans_39__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_3__dout),
    .if_empty_n(fifo_B_pe_Sextans_3__empty_n),
    .if_read(fifo_B_pe_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_3__din),
    .if_full_n(fifo_B_pe_Sextans_3__full_n),
    .if_write(fifo_B_pe_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_40
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_40__dout),
    .if_empty_n(fifo_B_pe_Sextans_40__empty_n),
    .if_read(fifo_B_pe_Sextans_40__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_40__din),
    .if_full_n(fifo_B_pe_Sextans_40__full_n),
    .if_write(fifo_B_pe_Sextans_40__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_41
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_41__dout),
    .if_empty_n(fifo_B_pe_Sextans_41__empty_n),
    .if_read(fifo_B_pe_Sextans_41__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_41__din),
    .if_full_n(fifo_B_pe_Sextans_41__full_n),
    .if_write(fifo_B_pe_Sextans_41__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_42
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_42__dout),
    .if_empty_n(fifo_B_pe_Sextans_42__empty_n),
    .if_read(fifo_B_pe_Sextans_42__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_42__din),
    .if_full_n(fifo_B_pe_Sextans_42__full_n),
    .if_write(fifo_B_pe_Sextans_42__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_43
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_43__dout),
    .if_empty_n(fifo_B_pe_Sextans_43__empty_n),
    .if_read(fifo_B_pe_Sextans_43__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_43__din),
    .if_full_n(fifo_B_pe_Sextans_43__full_n),
    .if_write(fifo_B_pe_Sextans_43__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_44
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_44__dout),
    .if_empty_n(fifo_B_pe_Sextans_44__empty_n),
    .if_read(fifo_B_pe_Sextans_44__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_44__din),
    .if_full_n(fifo_B_pe_Sextans_44__full_n),
    .if_write(fifo_B_pe_Sextans_44__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_45
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_45__dout),
    .if_empty_n(fifo_B_pe_Sextans_45__empty_n),
    .if_read(fifo_B_pe_Sextans_45__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_45__din),
    .if_full_n(fifo_B_pe_Sextans_45__full_n),
    .if_write(fifo_B_pe_Sextans_45__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_46
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_46__dout),
    .if_empty_n(fifo_B_pe_Sextans_46__empty_n),
    .if_read(fifo_B_pe_Sextans_46__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_46__din),
    .if_full_n(fifo_B_pe_Sextans_46__full_n),
    .if_write(fifo_B_pe_Sextans_46__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_47
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_47__dout),
    .if_empty_n(fifo_B_pe_Sextans_47__empty_n),
    .if_read(fifo_B_pe_Sextans_47__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_47__din),
    .if_full_n(fifo_B_pe_Sextans_47__full_n),
    .if_write(fifo_B_pe_Sextans_47__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_48
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_48__dout),
    .if_empty_n(fifo_B_pe_Sextans_48__empty_n),
    .if_read(fifo_B_pe_Sextans_48__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_48__din),
    .if_full_n(fifo_B_pe_Sextans_48__full_n),
    .if_write(fifo_B_pe_Sextans_48__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_49
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_49__dout),
    .if_empty_n(fifo_B_pe_Sextans_49__empty_n),
    .if_read(fifo_B_pe_Sextans_49__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_49__din),
    .if_full_n(fifo_B_pe_Sextans_49__full_n),
    .if_write(fifo_B_pe_Sextans_49__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_4__dout),
    .if_empty_n(fifo_B_pe_Sextans_4__empty_n),
    .if_read(fifo_B_pe_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_4__din),
    .if_full_n(fifo_B_pe_Sextans_4__full_n),
    .if_write(fifo_B_pe_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_50
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_50__dout),
    .if_empty_n(fifo_B_pe_Sextans_50__empty_n),
    .if_read(fifo_B_pe_Sextans_50__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_50__din),
    .if_full_n(fifo_B_pe_Sextans_50__full_n),
    .if_write(fifo_B_pe_Sextans_50__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_51
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_51__dout),
    .if_empty_n(fifo_B_pe_Sextans_51__empty_n),
    .if_read(fifo_B_pe_Sextans_51__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_51__din),
    .if_full_n(fifo_B_pe_Sextans_51__full_n),
    .if_write(fifo_B_pe_Sextans_51__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_52
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_52__dout),
    .if_empty_n(fifo_B_pe_Sextans_52__empty_n),
    .if_read(fifo_B_pe_Sextans_52__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_52__din),
    .if_full_n(fifo_B_pe_Sextans_52__full_n),
    .if_write(fifo_B_pe_Sextans_52__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_53
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_53__dout),
    .if_empty_n(fifo_B_pe_Sextans_53__empty_n),
    .if_read(fifo_B_pe_Sextans_53__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_53__din),
    .if_full_n(fifo_B_pe_Sextans_53__full_n),
    .if_write(fifo_B_pe_Sextans_53__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_54
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_54__dout),
    .if_empty_n(fifo_B_pe_Sextans_54__empty_n),
    .if_read(fifo_B_pe_Sextans_54__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_54__din),
    .if_full_n(fifo_B_pe_Sextans_54__full_n),
    .if_write(fifo_B_pe_Sextans_54__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_55
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_55__dout),
    .if_empty_n(fifo_B_pe_Sextans_55__empty_n),
    .if_read(fifo_B_pe_Sextans_55__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_55__din),
    .if_full_n(fifo_B_pe_Sextans_55__full_n),
    .if_write(fifo_B_pe_Sextans_55__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_56
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_56__dout),
    .if_empty_n(fifo_B_pe_Sextans_56__empty_n),
    .if_read(fifo_B_pe_Sextans_56__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_56__din),
    .if_full_n(fifo_B_pe_Sextans_56__full_n),
    .if_write(fifo_B_pe_Sextans_56__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_57
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_57__dout),
    .if_empty_n(fifo_B_pe_Sextans_57__empty_n),
    .if_read(fifo_B_pe_Sextans_57__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_57__din),
    .if_full_n(fifo_B_pe_Sextans_57__full_n),
    .if_write(fifo_B_pe_Sextans_57__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_58
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_58__dout),
    .if_empty_n(fifo_B_pe_Sextans_58__empty_n),
    .if_read(fifo_B_pe_Sextans_58__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_58__din),
    .if_full_n(fifo_B_pe_Sextans_58__full_n),
    .if_write(fifo_B_pe_Sextans_58__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_59
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_59__dout),
    .if_empty_n(fifo_B_pe_Sextans_59__empty_n),
    .if_read(fifo_B_pe_Sextans_59__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_59__din),
    .if_full_n(fifo_B_pe_Sextans_59__full_n),
    .if_write(fifo_B_pe_Sextans_59__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_5__dout),
    .if_empty_n(fifo_B_pe_Sextans_5__empty_n),
    .if_read(fifo_B_pe_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_5__din),
    .if_full_n(fifo_B_pe_Sextans_5__full_n),
    .if_write(fifo_B_pe_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_60
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_60__dout),
    .if_empty_n(fifo_B_pe_Sextans_60__empty_n),
    .if_read(fifo_B_pe_Sextans_60__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_60__din),
    .if_full_n(fifo_B_pe_Sextans_60__full_n),
    .if_write(fifo_B_pe_Sextans_60__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_61
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_61__dout),
    .if_empty_n(fifo_B_pe_Sextans_61__empty_n),
    .if_read(fifo_B_pe_Sextans_61__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_61__din),
    .if_full_n(fifo_B_pe_Sextans_61__full_n),
    .if_write(fifo_B_pe_Sextans_61__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_62
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_62__dout),
    .if_empty_n(fifo_B_pe_Sextans_62__empty_n),
    .if_read(fifo_B_pe_Sextans_62__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_62__din),
    .if_full_n(fifo_B_pe_Sextans_62__full_n),
    .if_write(fifo_B_pe_Sextans_62__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_63
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_63__dout),
    .if_empty_n(fifo_B_pe_Sextans_63__empty_n),
    .if_read(fifo_B_pe_Sextans_63__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_63__din),
    .if_full_n(fifo_B_pe_Sextans_63__full_n),
    .if_write(fifo_B_pe_Sextans_63__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_64
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_64__dout),
    .if_empty_n(fifo_B_pe_Sextans_64__empty_n),
    .if_read(fifo_B_pe_Sextans_64__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_64__din),
    .if_full_n(fifo_B_pe_Sextans_64__full_n),
    .if_write(fifo_B_pe_Sextans_64__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_65
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_65__dout),
    .if_empty_n(fifo_B_pe_Sextans_65__empty_n),
    .if_read(fifo_B_pe_Sextans_65__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_65__din),
    .if_full_n(fifo_B_pe_Sextans_65__full_n),
    .if_write(fifo_B_pe_Sextans_65__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_66
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_66__dout),
    .if_empty_n(fifo_B_pe_Sextans_66__empty_n),
    .if_read(fifo_B_pe_Sextans_66__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_66__din),
    .if_full_n(fifo_B_pe_Sextans_66__full_n),
    .if_write(fifo_B_pe_Sextans_66__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_67
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_67__dout),
    .if_empty_n(fifo_B_pe_Sextans_67__empty_n),
    .if_read(fifo_B_pe_Sextans_67__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_67__din),
    .if_full_n(fifo_B_pe_Sextans_67__full_n),
    .if_write(fifo_B_pe_Sextans_67__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_6__dout),
    .if_empty_n(fifo_B_pe_Sextans_6__empty_n),
    .if_read(fifo_B_pe_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_6__din),
    .if_full_n(fifo_B_pe_Sextans_6__full_n),
    .if_write(fifo_B_pe_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_7__dout),
    .if_empty_n(fifo_B_pe_Sextans_7__empty_n),
    .if_read(fifo_B_pe_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_7__din),
    .if_full_n(fifo_B_pe_Sextans_7__full_n),
    .if_write(fifo_B_pe_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_8__dout),
    .if_empty_n(fifo_B_pe_Sextans_8__empty_n),
    .if_read(fifo_B_pe_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_8__din),
    .if_full_n(fifo_B_pe_Sextans_8__full_n),
    .if_write(fifo_B_pe_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_pe_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_pe_Sextans_9__dout),
    .if_empty_n(fifo_B_pe_Sextans_9__empty_n),
    .if_read(fifo_B_pe_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_pe_Sextans_9__din),
    .if_full_n(fifo_B_pe_Sextans_9__full_n),
    .if_write(fifo_B_pe_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_0__dout),
    .if_empty_n(fifo_C_ch_Sextans_0__empty_n),
    .if_read(fifo_C_ch_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_0__din),
    .if_full_n(fifo_C_ch_Sextans_0__full_n),
    .if_write(fifo_C_ch_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_1__dout),
    .if_empty_n(fifo_C_ch_Sextans_1__empty_n),
    .if_read(fifo_C_ch_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_1__din),
    .if_full_n(fifo_C_ch_Sextans_1__full_n),
    .if_write(fifo_C_ch_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_2__dout),
    .if_empty_n(fifo_C_ch_Sextans_2__empty_n),
    .if_read(fifo_C_ch_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_2__din),
    .if_full_n(fifo_C_ch_Sextans_2__full_n),
    .if_write(fifo_C_ch_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_3__dout),
    .if_empty_n(fifo_C_ch_Sextans_3__empty_n),
    .if_read(fifo_C_ch_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_3__din),
    .if_full_n(fifo_C_ch_Sextans_3__full_n),
    .if_write(fifo_C_ch_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_4__dout),
    .if_empty_n(fifo_C_ch_Sextans_4__empty_n),
    .if_read(fifo_C_ch_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_4__din),
    .if_full_n(fifo_C_ch_Sextans_4__full_n),
    .if_write(fifo_C_ch_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_5__dout),
    .if_empty_n(fifo_C_ch_Sextans_5__empty_n),
    .if_read(fifo_C_ch_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_5__din),
    .if_full_n(fifo_C_ch_Sextans_5__full_n),
    .if_write(fifo_C_ch_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_6__dout),
    .if_empty_n(fifo_C_ch_Sextans_6__empty_n),
    .if_read(fifo_C_ch_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_6__din),
    .if_full_n(fifo_C_ch_Sextans_6__full_n),
    .if_write(fifo_C_ch_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_Sextans_7__dout),
    .if_empty_n(fifo_C_ch_Sextans_7__empty_n),
    .if_read(fifo_C_ch_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_Sextans_7__din),
    .if_full_n(fifo_C_ch_Sextans_7__full_n),
    .if_write(fifo_C_ch_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_0__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_0__empty_n),
    .if_read(fifo_C_ch_result_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_0__din),
    .if_full_n(fifo_C_ch_result_Sextans_0__full_n),
    .if_write(fifo_C_ch_result_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_1__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_1__empty_n),
    .if_read(fifo_C_ch_result_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_1__din),
    .if_full_n(fifo_C_ch_result_Sextans_1__full_n),
    .if_write(fifo_C_ch_result_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_2__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_2__empty_n),
    .if_read(fifo_C_ch_result_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_2__din),
    .if_full_n(fifo_C_ch_result_Sextans_2__full_n),
    .if_write(fifo_C_ch_result_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_3__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_3__empty_n),
    .if_read(fifo_C_ch_result_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_3__din),
    .if_full_n(fifo_C_ch_result_Sextans_3__full_n),
    .if_write(fifo_C_ch_result_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_4__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_4__empty_n),
    .if_read(fifo_C_ch_result_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_4__din),
    .if_full_n(fifo_C_ch_result_Sextans_4__full_n),
    .if_write(fifo_C_ch_result_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_5__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_5__empty_n),
    .if_read(fifo_C_ch_result_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_5__din),
    .if_full_n(fifo_C_ch_result_Sextans_5__full_n),
    .if_write(fifo_C_ch_result_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_6__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_6__empty_n),
    .if_read(fifo_C_ch_result_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_6__din),
    .if_full_n(fifo_C_ch_result_Sextans_6__full_n),
    .if_write(fifo_C_ch_result_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_Sextans_7__dout),
    .if_empty_n(fifo_C_ch_result_Sextans_7__empty_n),
    .if_read(fifo_C_ch_result_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_Sextans_7__din),
    .if_full_n(fifo_C_ch_result_Sextans_7__full_n),
    .if_write(fifo_C_ch_result_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_0__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_0__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_0__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_0__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_1__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_1__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_1__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_1__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_2__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_2__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_2__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_2__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_3__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_3__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_3__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_3__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_4__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_4__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_4__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_4__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_5__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_5__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_5__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_5__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_6__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_6__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_6__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_6__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_ch_result_alpha_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_ch_result_alpha_Sextans_7__dout),
    .if_empty_n(fifo_C_ch_result_alpha_Sextans_7__empty_n),
    .if_read(fifo_C_ch_result_alpha_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_ch_result_alpha_Sextans_7__din),
    .if_full_n(fifo_C_ch_result_alpha_Sextans_7__full_n),
    .if_write(fifo_C_ch_result_alpha_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_0__dout),
    .if_empty_n(fifo_C_pe_Sextans_0__empty_n),
    .if_read(fifo_C_pe_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_0__din),
    .if_full_n(fifo_C_pe_Sextans_0__full_n),
    .if_write(fifo_C_pe_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_10__dout),
    .if_empty_n(fifo_C_pe_Sextans_10__empty_n),
    .if_read(fifo_C_pe_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_10__din),
    .if_full_n(fifo_C_pe_Sextans_10__full_n),
    .if_write(fifo_C_pe_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_11__dout),
    .if_empty_n(fifo_C_pe_Sextans_11__empty_n),
    .if_read(fifo_C_pe_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_11__din),
    .if_full_n(fifo_C_pe_Sextans_11__full_n),
    .if_write(fifo_C_pe_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_12__dout),
    .if_empty_n(fifo_C_pe_Sextans_12__empty_n),
    .if_read(fifo_C_pe_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_12__din),
    .if_full_n(fifo_C_pe_Sextans_12__full_n),
    .if_write(fifo_C_pe_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_13__dout),
    .if_empty_n(fifo_C_pe_Sextans_13__empty_n),
    .if_read(fifo_C_pe_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_13__din),
    .if_full_n(fifo_C_pe_Sextans_13__full_n),
    .if_write(fifo_C_pe_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_14__dout),
    .if_empty_n(fifo_C_pe_Sextans_14__empty_n),
    .if_read(fifo_C_pe_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_14__din),
    .if_full_n(fifo_C_pe_Sextans_14__full_n),
    .if_write(fifo_C_pe_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_15__dout),
    .if_empty_n(fifo_C_pe_Sextans_15__empty_n),
    .if_read(fifo_C_pe_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_15__din),
    .if_full_n(fifo_C_pe_Sextans_15__full_n),
    .if_write(fifo_C_pe_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_1__dout),
    .if_empty_n(fifo_C_pe_Sextans_1__empty_n),
    .if_read(fifo_C_pe_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_1__din),
    .if_full_n(fifo_C_pe_Sextans_1__full_n),
    .if_write(fifo_C_pe_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_2__dout),
    .if_empty_n(fifo_C_pe_Sextans_2__empty_n),
    .if_read(fifo_C_pe_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_2__din),
    .if_full_n(fifo_C_pe_Sextans_2__full_n),
    .if_write(fifo_C_pe_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_3__dout),
    .if_empty_n(fifo_C_pe_Sextans_3__empty_n),
    .if_read(fifo_C_pe_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_3__din),
    .if_full_n(fifo_C_pe_Sextans_3__full_n),
    .if_write(fifo_C_pe_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_4__dout),
    .if_empty_n(fifo_C_pe_Sextans_4__empty_n),
    .if_read(fifo_C_pe_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_4__din),
    .if_full_n(fifo_C_pe_Sextans_4__full_n),
    .if_write(fifo_C_pe_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_5__dout),
    .if_empty_n(fifo_C_pe_Sextans_5__empty_n),
    .if_read(fifo_C_pe_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_5__din),
    .if_full_n(fifo_C_pe_Sextans_5__full_n),
    .if_write(fifo_C_pe_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_6__dout),
    .if_empty_n(fifo_C_pe_Sextans_6__empty_n),
    .if_read(fifo_C_pe_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_6__din),
    .if_full_n(fifo_C_pe_Sextans_6__full_n),
    .if_write(fifo_C_pe_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_7__dout),
    .if_empty_n(fifo_C_pe_Sextans_7__empty_n),
    .if_read(fifo_C_pe_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_7__din),
    .if_full_n(fifo_C_pe_Sextans_7__full_n),
    .if_write(fifo_C_pe_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_8__dout),
    .if_empty_n(fifo_C_pe_Sextans_8__empty_n),
    .if_read(fifo_C_pe_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_8__din),
    .if_full_n(fifo_C_pe_Sextans_8__full_n),
    .if_write(fifo_C_pe_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(257),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_pe_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_pe_Sextans_9__dout),
    .if_empty_n(fifo_C_pe_Sextans_9__empty_n),
    .if_read(fifo_C_pe_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_pe_Sextans_9__din),
    .if_full_n(fifo_C_pe_Sextans_9__full_n),
    .if_write(fifo_C_pe_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_0__dout),
    .if_empty_n(fifo_C_read_in_Sextans_0__empty_n),
    .if_read(fifo_C_read_in_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_0__din),
    .if_full_n(fifo_C_read_in_Sextans_0__full_n),
    .if_write(fifo_C_read_in_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_1__dout),
    .if_empty_n(fifo_C_read_in_Sextans_1__empty_n),
    .if_read(fifo_C_read_in_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_1__din),
    .if_full_n(fifo_C_read_in_Sextans_1__full_n),
    .if_write(fifo_C_read_in_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_2__dout),
    .if_empty_n(fifo_C_read_in_Sextans_2__empty_n),
    .if_read(fifo_C_read_in_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_2__din),
    .if_full_n(fifo_C_read_in_Sextans_2__full_n),
    .if_write(fifo_C_read_in_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_3__dout),
    .if_empty_n(fifo_C_read_in_Sextans_3__empty_n),
    .if_read(fifo_C_read_in_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_3__din),
    .if_full_n(fifo_C_read_in_Sextans_3__full_n),
    .if_write(fifo_C_read_in_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_4__dout),
    .if_empty_n(fifo_C_read_in_Sextans_4__empty_n),
    .if_read(fifo_C_read_in_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_4__din),
    .if_full_n(fifo_C_read_in_Sextans_4__full_n),
    .if_write(fifo_C_read_in_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_5__dout),
    .if_empty_n(fifo_C_read_in_Sextans_5__empty_n),
    .if_read(fifo_C_read_in_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_5__din),
    .if_full_n(fifo_C_read_in_Sextans_5__full_n),
    .if_write(fifo_C_read_in_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_6__dout),
    .if_empty_n(fifo_C_read_in_Sextans_6__empty_n),
    .if_read(fifo_C_read_in_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_6__din),
    .if_full_n(fifo_C_read_in_Sextans_6__full_n),
    .if_write(fifo_C_read_in_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_Sextans_7__dout),
    .if_empty_n(fifo_C_read_in_Sextans_7__empty_n),
    .if_read(fifo_C_read_in_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_Sextans_7__din),
    .if_full_n(fifo_C_read_in_Sextans_7__full_n),
    .if_write(fifo_C_read_in_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_0__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_0__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_0__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_0__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_1__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_1__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_1__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_1__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_2__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_2__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_2__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_2__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_3__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_3__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_3__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_3__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_4__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_4__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_4__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_4__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_5__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_5__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_5__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_5__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_6__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_6__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_6__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_6__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_read_in_beta_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_read_in_beta_Sextans_7__dout),
    .if_empty_n(fifo_C_read_in_beta_Sextans_7__empty_n),
    .if_read(fifo_C_read_in_beta_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_read_in_beta_Sextans_7__din),
    .if_full_n(fifo_C_read_in_beta_Sextans_7__full_n),
    .if_write(fifo_C_read_in_beta_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_0__dout),
    .if_empty_n(fifo_aBvec_Sextans_0__empty_n),
    .if_read(fifo_aBvec_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_0__din),
    .if_full_n(fifo_aBvec_Sextans_0__full_n),
    .if_write(fifo_aBvec_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_10__dout),
    .if_empty_n(fifo_aBvec_Sextans_10__empty_n),
    .if_read(fifo_aBvec_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_10__din),
    .if_full_n(fifo_aBvec_Sextans_10__full_n),
    .if_write(fifo_aBvec_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_11__dout),
    .if_empty_n(fifo_aBvec_Sextans_11__empty_n),
    .if_read(fifo_aBvec_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_11__din),
    .if_full_n(fifo_aBvec_Sextans_11__full_n),
    .if_write(fifo_aBvec_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_12__dout),
    .if_empty_n(fifo_aBvec_Sextans_12__empty_n),
    .if_read(fifo_aBvec_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_12__din),
    .if_full_n(fifo_aBvec_Sextans_12__full_n),
    .if_write(fifo_aBvec_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_13__dout),
    .if_empty_n(fifo_aBvec_Sextans_13__empty_n),
    .if_read(fifo_aBvec_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_13__din),
    .if_full_n(fifo_aBvec_Sextans_13__full_n),
    .if_write(fifo_aBvec_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_14__dout),
    .if_empty_n(fifo_aBvec_Sextans_14__empty_n),
    .if_read(fifo_aBvec_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_14__din),
    .if_full_n(fifo_aBvec_Sextans_14__full_n),
    .if_write(fifo_aBvec_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_15__dout),
    .if_empty_n(fifo_aBvec_Sextans_15__empty_n),
    .if_read(fifo_aBvec_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_15__din),
    .if_full_n(fifo_aBvec_Sextans_15__full_n),
    .if_write(fifo_aBvec_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_16__dout),
    .if_empty_n(fifo_aBvec_Sextans_16__empty_n),
    .if_read(fifo_aBvec_Sextans_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_16__din),
    .if_full_n(fifo_aBvec_Sextans_16__full_n),
    .if_write(fifo_aBvec_Sextans_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_17__dout),
    .if_empty_n(fifo_aBvec_Sextans_17__empty_n),
    .if_read(fifo_aBvec_Sextans_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_17__din),
    .if_full_n(fifo_aBvec_Sextans_17__full_n),
    .if_write(fifo_aBvec_Sextans_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_18
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_18__dout),
    .if_empty_n(fifo_aBvec_Sextans_18__empty_n),
    .if_read(fifo_aBvec_Sextans_18__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_18__din),
    .if_full_n(fifo_aBvec_Sextans_18__full_n),
    .if_write(fifo_aBvec_Sextans_18__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_19
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_19__dout),
    .if_empty_n(fifo_aBvec_Sextans_19__empty_n),
    .if_read(fifo_aBvec_Sextans_19__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_19__din),
    .if_full_n(fifo_aBvec_Sextans_19__full_n),
    .if_write(fifo_aBvec_Sextans_19__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_1__dout),
    .if_empty_n(fifo_aBvec_Sextans_1__empty_n),
    .if_read(fifo_aBvec_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_1__din),
    .if_full_n(fifo_aBvec_Sextans_1__full_n),
    .if_write(fifo_aBvec_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_20
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_20__dout),
    .if_empty_n(fifo_aBvec_Sextans_20__empty_n),
    .if_read(fifo_aBvec_Sextans_20__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_20__din),
    .if_full_n(fifo_aBvec_Sextans_20__full_n),
    .if_write(fifo_aBvec_Sextans_20__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_21
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_21__dout),
    .if_empty_n(fifo_aBvec_Sextans_21__empty_n),
    .if_read(fifo_aBvec_Sextans_21__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_21__din),
    .if_full_n(fifo_aBvec_Sextans_21__full_n),
    .if_write(fifo_aBvec_Sextans_21__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_22
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_22__dout),
    .if_empty_n(fifo_aBvec_Sextans_22__empty_n),
    .if_read(fifo_aBvec_Sextans_22__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_22__din),
    .if_full_n(fifo_aBvec_Sextans_22__full_n),
    .if_write(fifo_aBvec_Sextans_22__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_23
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_23__dout),
    .if_empty_n(fifo_aBvec_Sextans_23__empty_n),
    .if_read(fifo_aBvec_Sextans_23__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_23__din),
    .if_full_n(fifo_aBvec_Sextans_23__full_n),
    .if_write(fifo_aBvec_Sextans_23__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_24
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_24__dout),
    .if_empty_n(fifo_aBvec_Sextans_24__empty_n),
    .if_read(fifo_aBvec_Sextans_24__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_24__din),
    .if_full_n(fifo_aBvec_Sextans_24__full_n),
    .if_write(fifo_aBvec_Sextans_24__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_25
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_25__dout),
    .if_empty_n(fifo_aBvec_Sextans_25__empty_n),
    .if_read(fifo_aBvec_Sextans_25__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_25__din),
    .if_full_n(fifo_aBvec_Sextans_25__full_n),
    .if_write(fifo_aBvec_Sextans_25__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_26
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_26__dout),
    .if_empty_n(fifo_aBvec_Sextans_26__empty_n),
    .if_read(fifo_aBvec_Sextans_26__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_26__din),
    .if_full_n(fifo_aBvec_Sextans_26__full_n),
    .if_write(fifo_aBvec_Sextans_26__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_27
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_27__dout),
    .if_empty_n(fifo_aBvec_Sextans_27__empty_n),
    .if_read(fifo_aBvec_Sextans_27__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_27__din),
    .if_full_n(fifo_aBvec_Sextans_27__full_n),
    .if_write(fifo_aBvec_Sextans_27__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_28
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_28__dout),
    .if_empty_n(fifo_aBvec_Sextans_28__empty_n),
    .if_read(fifo_aBvec_Sextans_28__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_28__din),
    .if_full_n(fifo_aBvec_Sextans_28__full_n),
    .if_write(fifo_aBvec_Sextans_28__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_29
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_29__dout),
    .if_empty_n(fifo_aBvec_Sextans_29__empty_n),
    .if_read(fifo_aBvec_Sextans_29__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_29__din),
    .if_full_n(fifo_aBvec_Sextans_29__full_n),
    .if_write(fifo_aBvec_Sextans_29__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_2__dout),
    .if_empty_n(fifo_aBvec_Sextans_2__empty_n),
    .if_read(fifo_aBvec_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_2__din),
    .if_full_n(fifo_aBvec_Sextans_2__full_n),
    .if_write(fifo_aBvec_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_30
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_30__dout),
    .if_empty_n(fifo_aBvec_Sextans_30__empty_n),
    .if_read(fifo_aBvec_Sextans_30__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_30__din),
    .if_full_n(fifo_aBvec_Sextans_30__full_n),
    .if_write(fifo_aBvec_Sextans_30__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_31
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_31__dout),
    .if_empty_n(fifo_aBvec_Sextans_31__empty_n),
    .if_read(fifo_aBvec_Sextans_31__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_31__din),
    .if_full_n(fifo_aBvec_Sextans_31__full_n),
    .if_write(fifo_aBvec_Sextans_31__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_32
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_32__dout),
    .if_empty_n(fifo_aBvec_Sextans_32__empty_n),
    .if_read(fifo_aBvec_Sextans_32__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_32__din),
    .if_full_n(fifo_aBvec_Sextans_32__full_n),
    .if_write(fifo_aBvec_Sextans_32__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_33
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_33__dout),
    .if_empty_n(fifo_aBvec_Sextans_33__empty_n),
    .if_read(fifo_aBvec_Sextans_33__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_33__din),
    .if_full_n(fifo_aBvec_Sextans_33__full_n),
    .if_write(fifo_aBvec_Sextans_33__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_34
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_34__dout),
    .if_empty_n(fifo_aBvec_Sextans_34__empty_n),
    .if_read(fifo_aBvec_Sextans_34__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_34__din),
    .if_full_n(fifo_aBvec_Sextans_34__full_n),
    .if_write(fifo_aBvec_Sextans_34__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_35
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_35__dout),
    .if_empty_n(fifo_aBvec_Sextans_35__empty_n),
    .if_read(fifo_aBvec_Sextans_35__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_35__din),
    .if_full_n(fifo_aBvec_Sextans_35__full_n),
    .if_write(fifo_aBvec_Sextans_35__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_36
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_36__dout),
    .if_empty_n(fifo_aBvec_Sextans_36__empty_n),
    .if_read(fifo_aBvec_Sextans_36__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_36__din),
    .if_full_n(fifo_aBvec_Sextans_36__full_n),
    .if_write(fifo_aBvec_Sextans_36__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_37
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_37__dout),
    .if_empty_n(fifo_aBvec_Sextans_37__empty_n),
    .if_read(fifo_aBvec_Sextans_37__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_37__din),
    .if_full_n(fifo_aBvec_Sextans_37__full_n),
    .if_write(fifo_aBvec_Sextans_37__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_38
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_38__dout),
    .if_empty_n(fifo_aBvec_Sextans_38__empty_n),
    .if_read(fifo_aBvec_Sextans_38__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_38__din),
    .if_full_n(fifo_aBvec_Sextans_38__full_n),
    .if_write(fifo_aBvec_Sextans_38__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_39
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_39__dout),
    .if_empty_n(fifo_aBvec_Sextans_39__empty_n),
    .if_read(fifo_aBvec_Sextans_39__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_39__din),
    .if_full_n(fifo_aBvec_Sextans_39__full_n),
    .if_write(fifo_aBvec_Sextans_39__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_3__dout),
    .if_empty_n(fifo_aBvec_Sextans_3__empty_n),
    .if_read(fifo_aBvec_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_3__din),
    .if_full_n(fifo_aBvec_Sextans_3__full_n),
    .if_write(fifo_aBvec_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_40
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_40__dout),
    .if_empty_n(fifo_aBvec_Sextans_40__empty_n),
    .if_read(fifo_aBvec_Sextans_40__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_40__din),
    .if_full_n(fifo_aBvec_Sextans_40__full_n),
    .if_write(fifo_aBvec_Sextans_40__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_41
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_41__dout),
    .if_empty_n(fifo_aBvec_Sextans_41__empty_n),
    .if_read(fifo_aBvec_Sextans_41__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_41__din),
    .if_full_n(fifo_aBvec_Sextans_41__full_n),
    .if_write(fifo_aBvec_Sextans_41__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_42
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_42__dout),
    .if_empty_n(fifo_aBvec_Sextans_42__empty_n),
    .if_read(fifo_aBvec_Sextans_42__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_42__din),
    .if_full_n(fifo_aBvec_Sextans_42__full_n),
    .if_write(fifo_aBvec_Sextans_42__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_43
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_43__dout),
    .if_empty_n(fifo_aBvec_Sextans_43__empty_n),
    .if_read(fifo_aBvec_Sextans_43__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_43__din),
    .if_full_n(fifo_aBvec_Sextans_43__full_n),
    .if_write(fifo_aBvec_Sextans_43__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_44
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_44__dout),
    .if_empty_n(fifo_aBvec_Sextans_44__empty_n),
    .if_read(fifo_aBvec_Sextans_44__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_44__din),
    .if_full_n(fifo_aBvec_Sextans_44__full_n),
    .if_write(fifo_aBvec_Sextans_44__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_45
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_45__dout),
    .if_empty_n(fifo_aBvec_Sextans_45__empty_n),
    .if_read(fifo_aBvec_Sextans_45__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_45__din),
    .if_full_n(fifo_aBvec_Sextans_45__full_n),
    .if_write(fifo_aBvec_Sextans_45__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_46
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_46__dout),
    .if_empty_n(fifo_aBvec_Sextans_46__empty_n),
    .if_read(fifo_aBvec_Sextans_46__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_46__din),
    .if_full_n(fifo_aBvec_Sextans_46__full_n),
    .if_write(fifo_aBvec_Sextans_46__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_47
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_47__dout),
    .if_empty_n(fifo_aBvec_Sextans_47__empty_n),
    .if_read(fifo_aBvec_Sextans_47__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_47__din),
    .if_full_n(fifo_aBvec_Sextans_47__full_n),
    .if_write(fifo_aBvec_Sextans_47__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_48
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_48__dout),
    .if_empty_n(fifo_aBvec_Sextans_48__empty_n),
    .if_read(fifo_aBvec_Sextans_48__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_48__din),
    .if_full_n(fifo_aBvec_Sextans_48__full_n),
    .if_write(fifo_aBvec_Sextans_48__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_49
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_49__dout),
    .if_empty_n(fifo_aBvec_Sextans_49__empty_n),
    .if_read(fifo_aBvec_Sextans_49__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_49__din),
    .if_full_n(fifo_aBvec_Sextans_49__full_n),
    .if_write(fifo_aBvec_Sextans_49__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_4__dout),
    .if_empty_n(fifo_aBvec_Sextans_4__empty_n),
    .if_read(fifo_aBvec_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_4__din),
    .if_full_n(fifo_aBvec_Sextans_4__full_n),
    .if_write(fifo_aBvec_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_50
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_50__dout),
    .if_empty_n(fifo_aBvec_Sextans_50__empty_n),
    .if_read(fifo_aBvec_Sextans_50__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_50__din),
    .if_full_n(fifo_aBvec_Sextans_50__full_n),
    .if_write(fifo_aBvec_Sextans_50__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_51
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_51__dout),
    .if_empty_n(fifo_aBvec_Sextans_51__empty_n),
    .if_read(fifo_aBvec_Sextans_51__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_51__din),
    .if_full_n(fifo_aBvec_Sextans_51__full_n),
    .if_write(fifo_aBvec_Sextans_51__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_52
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_52__dout),
    .if_empty_n(fifo_aBvec_Sextans_52__empty_n),
    .if_read(fifo_aBvec_Sextans_52__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_52__din),
    .if_full_n(fifo_aBvec_Sextans_52__full_n),
    .if_write(fifo_aBvec_Sextans_52__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_53
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_53__dout),
    .if_empty_n(fifo_aBvec_Sextans_53__empty_n),
    .if_read(fifo_aBvec_Sextans_53__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_53__din),
    .if_full_n(fifo_aBvec_Sextans_53__full_n),
    .if_write(fifo_aBvec_Sextans_53__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_54
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_54__dout),
    .if_empty_n(fifo_aBvec_Sextans_54__empty_n),
    .if_read(fifo_aBvec_Sextans_54__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_54__din),
    .if_full_n(fifo_aBvec_Sextans_54__full_n),
    .if_write(fifo_aBvec_Sextans_54__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_55
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_55__dout),
    .if_empty_n(fifo_aBvec_Sextans_55__empty_n),
    .if_read(fifo_aBvec_Sextans_55__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_55__din),
    .if_full_n(fifo_aBvec_Sextans_55__full_n),
    .if_write(fifo_aBvec_Sextans_55__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_56
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_56__dout),
    .if_empty_n(fifo_aBvec_Sextans_56__empty_n),
    .if_read(fifo_aBvec_Sextans_56__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_56__din),
    .if_full_n(fifo_aBvec_Sextans_56__full_n),
    .if_write(fifo_aBvec_Sextans_56__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_57
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_57__dout),
    .if_empty_n(fifo_aBvec_Sextans_57__empty_n),
    .if_read(fifo_aBvec_Sextans_57__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_57__din),
    .if_full_n(fifo_aBvec_Sextans_57__full_n),
    .if_write(fifo_aBvec_Sextans_57__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_58
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_58__dout),
    .if_empty_n(fifo_aBvec_Sextans_58__empty_n),
    .if_read(fifo_aBvec_Sextans_58__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_58__din),
    .if_full_n(fifo_aBvec_Sextans_58__full_n),
    .if_write(fifo_aBvec_Sextans_58__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_59
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_59__dout),
    .if_empty_n(fifo_aBvec_Sextans_59__empty_n),
    .if_read(fifo_aBvec_Sextans_59__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_59__din),
    .if_full_n(fifo_aBvec_Sextans_59__full_n),
    .if_write(fifo_aBvec_Sextans_59__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_5__dout),
    .if_empty_n(fifo_aBvec_Sextans_5__empty_n),
    .if_read(fifo_aBvec_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_5__din),
    .if_full_n(fifo_aBvec_Sextans_5__full_n),
    .if_write(fifo_aBvec_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_60
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_60__dout),
    .if_empty_n(fifo_aBvec_Sextans_60__empty_n),
    .if_read(fifo_aBvec_Sextans_60__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_60__din),
    .if_full_n(fifo_aBvec_Sextans_60__full_n),
    .if_write(fifo_aBvec_Sextans_60__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_61
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_61__dout),
    .if_empty_n(fifo_aBvec_Sextans_61__empty_n),
    .if_read(fifo_aBvec_Sextans_61__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_61__din),
    .if_full_n(fifo_aBvec_Sextans_61__full_n),
    .if_write(fifo_aBvec_Sextans_61__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_62
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_62__dout),
    .if_empty_n(fifo_aBvec_Sextans_62__empty_n),
    .if_read(fifo_aBvec_Sextans_62__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_62__din),
    .if_full_n(fifo_aBvec_Sextans_62__full_n),
    .if_write(fifo_aBvec_Sextans_62__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_63
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_63__dout),
    .if_empty_n(fifo_aBvec_Sextans_63__empty_n),
    .if_read(fifo_aBvec_Sextans_63__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_63__din),
    .if_full_n(fifo_aBvec_Sextans_63__full_n),
    .if_write(fifo_aBvec_Sextans_63__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_6__dout),
    .if_empty_n(fifo_aBvec_Sextans_6__empty_n),
    .if_read(fifo_aBvec_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_6__din),
    .if_full_n(fifo_aBvec_Sextans_6__full_n),
    .if_write(fifo_aBvec_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_7__dout),
    .if_empty_n(fifo_aBvec_Sextans_7__empty_n),
    .if_read(fifo_aBvec_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_7__din),
    .if_full_n(fifo_aBvec_Sextans_7__full_n),
    .if_write(fifo_aBvec_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_8__dout),
    .if_empty_n(fifo_aBvec_Sextans_8__empty_n),
    .if_read(fifo_aBvec_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_8__din),
    .if_full_n(fifo_aBvec_Sextans_8__full_n),
    .if_write(fifo_aBvec_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(275),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_aBvec_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_aBvec_Sextans_9__dout),
    .if_empty_n(fifo_aBvec_Sextans_9__empty_n),
    .if_read(fifo_aBvec_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_aBvec_Sextans_9__din),
    .if_full_n(fifo_aBvec_Sextans_9__full_n),
    .if_write(fifo_aBvec_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_0__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_0__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_0__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_0__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_10__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_10__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_10__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_10__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_11__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_11__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_11__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_11__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_12__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_12__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_12__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_12__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_13__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_13__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_13__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_13__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_14__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_14__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_14__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_14__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_15__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_15__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_15__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_15__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_16__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_16__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_16__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_16__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_1__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_1__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_1__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_1__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_2__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_2__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_2__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_2__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_3__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_3__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_3__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_3__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_4__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_4__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_4__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_4__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_5__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_5__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_5__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_5__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_6__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_6__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_6__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_6__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_7__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_7__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_7__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_7__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_8__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_8__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_8__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_8__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_Sextans_9__dout),
    .if_empty_n(fifo_edge_list_ptr_Sextans_9__empty_n),
    .if_read(fifo_edge_list_ptr_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_Sextans_9__din),
    .if_full_n(fifo_edge_list_ptr_Sextans_9__full_n),
    .if_write(fifo_edge_list_ptr_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_0__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_0__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_0__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_0__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_10__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_10__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_10__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_10__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_11__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_11__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_11__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_11__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_12__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_12__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_12__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_12__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_13__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_13__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_13__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_13__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_14__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_14__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_14__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_14__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_15__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_15__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_15__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_15__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_1__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_1__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_1__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_1__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_2__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_2__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_2__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_2__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_3__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_3__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_3__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_3__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_4__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_4__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_4__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_4__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_5__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_5__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_5__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_5__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_6__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_6__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_6__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_6__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_7__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_7__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_7__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_7__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_8__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_8__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_8__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_8__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_edge_list_ptr_to_Cmtx_Sextans_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_9__dout),
    .if_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_9__empty_n),
    .if_read(fifo_edge_list_ptr_to_Cmtx_Sextans_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_edge_list_ptr_to_Cmtx_Sextans_9__din),
    .if_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_9__full_n),
    .if_write(fifo_edge_list_ptr_to_Cmtx_Sextans_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_0__dout),
    .if_empty_n(wrC_inst_Sextans_0__empty_n),
    .if_read(wrC_inst_Sextans_0__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_0__din),
    .if_full_n(wrC_inst_Sextans_0__full_n),
    .if_write(wrC_inst_Sextans_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_1__dout),
    .if_empty_n(wrC_inst_Sextans_1__empty_n),
    .if_read(wrC_inst_Sextans_1__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_1__din),
    .if_full_n(wrC_inst_Sextans_1__full_n),
    .if_write(wrC_inst_Sextans_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_2__dout),
    .if_empty_n(wrC_inst_Sextans_2__empty_n),
    .if_read(wrC_inst_Sextans_2__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_2__din),
    .if_full_n(wrC_inst_Sextans_2__full_n),
    .if_write(wrC_inst_Sextans_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_3__dout),
    .if_empty_n(wrC_inst_Sextans_3__empty_n),
    .if_read(wrC_inst_Sextans_3__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_3__din),
    .if_full_n(wrC_inst_Sextans_3__full_n),
    .if_write(wrC_inst_Sextans_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_4__dout),
    .if_empty_n(wrC_inst_Sextans_4__empty_n),
    .if_read(wrC_inst_Sextans_4__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_4__din),
    .if_full_n(wrC_inst_Sextans_4__full_n),
    .if_write(wrC_inst_Sextans_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_5__dout),
    .if_empty_n(wrC_inst_Sextans_5__empty_n),
    .if_read(wrC_inst_Sextans_5__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_5__din),
    .if_full_n(wrC_inst_Sextans_5__full_n),
    .if_write(wrC_inst_Sextans_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_6__dout),
    .if_empty_n(wrC_inst_Sextans_6__empty_n),
    .if_read(wrC_inst_Sextans_6__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_6__din),
    .if_full_n(wrC_inst_Sextans_6__full_n),
    .if_write(wrC_inst_Sextans_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  wrC_inst_Sextans_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(wrC_inst_Sextans_7__dout),
    .if_empty_n(wrC_inst_Sextans_7__empty_n),
    .if_read(wrC_inst_Sextans_7__read),
    .if_read_ce(1'b1),
    .if_din(wrC_inst_Sextans_7__din),
    .if_full_n(wrC_inst_Sextans_7__full_n),
    .if_write(wrC_inst_Sextans_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_0__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_0__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_0__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_0__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_0__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_0__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_0__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_0__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_0__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_0__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_0__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_0__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_0__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_1__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_1__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_1__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_1__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_1__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_1__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_1__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_1__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_1__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_1__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_1__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_1__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_1__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_2__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_2__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_2__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_2__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_2__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_2__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_2__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_2__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_2__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_2__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_2__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_2__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_2__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_2__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_3__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_3__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_3__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_3__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_3__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_3__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_3__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_3__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_3__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_3__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_3__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_3__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_3__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_3__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_4__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_4__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_4__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_4__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_4__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_4__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_4__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_4__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_4__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_4__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_4__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_4__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_4__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_4__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_5__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_5__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_5__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_5__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_5__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_5__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_5__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_5__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_5__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_5__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_5__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_5__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_5__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_5__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_6__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_6__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_6__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_6__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_6__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_6__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_6__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_6__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_6__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_6__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_6__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_6__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_6__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_6__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvAddFloatv
  FloatvAddFloatv_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvAddFloatv_7__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_Sextans_7__din),
    .fifo_out_full_n(fifo_C_ch_Sextans_7__full_n),
    .fifo_out_write(fifo_C_ch_Sextans_7__write),
    .fifo_in0_s_dout(fifo_C_ch_result_alpha_Sextans_7__dout),
    .fifo_in0_peek_dout(fifo_C_ch_result_alpha_Sextans_7__dout),
    .fifo_in0_s_empty_n(fifo_C_ch_result_alpha_Sextans_7__empty_n),
    .fifo_in0_peek_empty_n(fifo_C_ch_result_alpha_Sextans_7__empty_n),
    .fifo_in0_s_read(fifo_C_ch_result_alpha_Sextans_7__read),
    .fifo_in0_peek_read(),
    .fifo_in1_s_dout(fifo_C_read_in_beta_Sextans_7__dout),
    .fifo_in1_peek_dout(fifo_C_read_in_beta_Sextans_7__dout),
    .fifo_in1_s_empty_n(fifo_C_read_in_beta_Sextans_7__empty_n),
    .fifo_in1_peek_empty_n(fifo_C_read_in_beta_Sextans_7__empty_n),
    .fifo_in1_s_read(fifo_C_read_in_beta_Sextans_7__read),
    .fifo_in1_peek_read()
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_0__ap_start),
    .ap_done(FloatvMultConst_0__ap_done),
    .ap_idle(FloatvMultConst_0__ap_idle),
    .ap_ready(FloatvMultConst_0__ap_ready),
    .M(FloatvMultConst_0___M__q0),
    .P_N(FloatvMultConst_0___P_N__q0),
    .alpha_u(FloatvMultConst_0___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_0__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_0__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_0__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_0__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_0__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_0__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_0__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_0__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_1__ap_start),
    .ap_done(FloatvMultConst_1__ap_done),
    .ap_idle(FloatvMultConst_1__ap_idle),
    .ap_ready(FloatvMultConst_1__ap_ready),
    .M(FloatvMultConst_1___M__q0),
    .P_N(FloatvMultConst_1___P_N__q0),
    .alpha_u(FloatvMultConst_1___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_1__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_1__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_1__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_1__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_1__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_1__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_1__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_1__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_2__ap_start),
    .ap_done(FloatvMultConst_2__ap_done),
    .ap_idle(FloatvMultConst_2__ap_idle),
    .ap_ready(FloatvMultConst_2__ap_ready),
    .M(FloatvMultConst_2___M__q0),
    .P_N(FloatvMultConst_2___P_N__q0),
    .alpha_u(FloatvMultConst_2___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_2__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_2__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_2__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_2__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_2__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_2__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_2__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_2__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_3__ap_start),
    .ap_done(FloatvMultConst_3__ap_done),
    .ap_idle(FloatvMultConst_3__ap_idle),
    .ap_ready(FloatvMultConst_3__ap_ready),
    .M(FloatvMultConst_3___M__q0),
    .P_N(FloatvMultConst_3___P_N__q0),
    .alpha_u(FloatvMultConst_3___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_3__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_3__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_3__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_3__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_3__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_3__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_3__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_3__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_4__ap_start),
    .ap_done(FloatvMultConst_4__ap_done),
    .ap_idle(FloatvMultConst_4__ap_idle),
    .ap_ready(FloatvMultConst_4__ap_ready),
    .M(FloatvMultConst_4___M__q0),
    .P_N(FloatvMultConst_4___P_N__q0),
    .alpha_u(FloatvMultConst_4___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_4__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_4__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_4__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_4__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_4__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_4__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_4__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_4__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_5__ap_start),
    .ap_done(FloatvMultConst_5__ap_done),
    .ap_idle(FloatvMultConst_5__ap_idle),
    .ap_ready(FloatvMultConst_5__ap_ready),
    .M(FloatvMultConst_5___M__q0),
    .P_N(FloatvMultConst_5___P_N__q0),
    .alpha_u(FloatvMultConst_5___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_5__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_5__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_5__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_5__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_5__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_5__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_5__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_5__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_6__ap_start),
    .ap_done(FloatvMultConst_6__ap_done),
    .ap_idle(FloatvMultConst_6__ap_idle),
    .ap_ready(FloatvMultConst_6__ap_ready),
    .M(FloatvMultConst_6___M__q0),
    .P_N(FloatvMultConst_6___P_N__q0),
    .alpha_u(FloatvMultConst_6___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_6__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_6__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_6__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_6__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_6__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_6__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_6__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_6__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_7__ap_start),
    .ap_done(FloatvMultConst_7__ap_done),
    .ap_idle(FloatvMultConst_7__ap_idle),
    .ap_ready(FloatvMultConst_7__ap_ready),
    .M(FloatvMultConst_7___M__q0),
    .P_N(FloatvMultConst_7___P_N__q0),
    .alpha_u(FloatvMultConst_7___beta_u__q0),
    .fifo_in_s_dout(fifo_C_read_in_Sextans_7__dout),
    .fifo_in_peek_dout(fifo_C_read_in_Sextans_7__dout),
    .fifo_in_s_empty_n(fifo_C_read_in_Sextans_7__empty_n),
    .fifo_in_peek_empty_n(fifo_C_read_in_Sextans_7__empty_n),
    .fifo_in_s_read(fifo_C_read_in_Sextans_7__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_read_in_beta_Sextans_7__din),
    .fifo_out_full_n(fifo_C_read_in_beta_Sextans_7__full_n),
    .fifo_out_write(fifo_C_read_in_beta_Sextans_7__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_8__ap_start),
    .ap_done(FloatvMultConst_8__ap_done),
    .ap_idle(FloatvMultConst_8__ap_idle),
    .ap_ready(FloatvMultConst_8__ap_ready),
    .M(FloatvMultConst_8___M__q0),
    .P_N(FloatvMultConst_8___P_N__q0),
    .alpha_u(FloatvMultConst_8___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_0__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_0__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_0__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_0__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_0__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_0__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_0__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_0__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_9__ap_start),
    .ap_done(FloatvMultConst_9__ap_done),
    .ap_idle(FloatvMultConst_9__ap_idle),
    .ap_ready(FloatvMultConst_9__ap_ready),
    .M(FloatvMultConst_9___M__q0),
    .P_N(FloatvMultConst_9___P_N__q0),
    .alpha_u(FloatvMultConst_9___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_1__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_1__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_1__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_1__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_1__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_1__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_1__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_1__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_10__ap_start),
    .ap_done(FloatvMultConst_10__ap_done),
    .ap_idle(FloatvMultConst_10__ap_idle),
    .ap_ready(FloatvMultConst_10__ap_ready),
    .M(FloatvMultConst_10___M__q0),
    .P_N(FloatvMultConst_10___P_N__q0),
    .alpha_u(FloatvMultConst_10___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_2__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_2__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_2__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_2__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_2__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_2__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_2__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_2__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_11__ap_start),
    .ap_done(FloatvMultConst_11__ap_done),
    .ap_idle(FloatvMultConst_11__ap_idle),
    .ap_ready(FloatvMultConst_11__ap_ready),
    .M(FloatvMultConst_11___M__q0),
    .P_N(FloatvMultConst_11___P_N__q0),
    .alpha_u(FloatvMultConst_11___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_3__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_3__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_3__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_3__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_3__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_3__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_3__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_3__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_12__ap_start),
    .ap_done(FloatvMultConst_12__ap_done),
    .ap_idle(FloatvMultConst_12__ap_idle),
    .ap_ready(FloatvMultConst_12__ap_ready),
    .M(FloatvMultConst_12___M__q0),
    .P_N(FloatvMultConst_12___P_N__q0),
    .alpha_u(FloatvMultConst_12___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_4__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_4__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_4__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_4__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_4__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_4__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_4__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_4__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_13__ap_start),
    .ap_done(FloatvMultConst_13__ap_done),
    .ap_idle(FloatvMultConst_13__ap_idle),
    .ap_ready(FloatvMultConst_13__ap_ready),
    .M(FloatvMultConst_13___M__q0),
    .P_N(FloatvMultConst_13___P_N__q0),
    .alpha_u(FloatvMultConst_13___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_5__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_5__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_5__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_5__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_5__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_5__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_5__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_5__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_14__ap_start),
    .ap_done(FloatvMultConst_14__ap_done),
    .ap_idle(FloatvMultConst_14__ap_idle),
    .ap_ready(FloatvMultConst_14__ap_ready),
    .M(FloatvMultConst_14___M__q0),
    .P_N(FloatvMultConst_14___P_N__q0),
    .alpha_u(FloatvMultConst_14___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_6__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_6__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_6__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_6__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_6__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_6__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_6__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_6__write)
  );


  (* keep_hierarchy = "yes" *) FloatvMultConst
  FloatvMultConst_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(FloatvMultConst_15__ap_start),
    .ap_done(FloatvMultConst_15__ap_done),
    .ap_idle(FloatvMultConst_15__ap_idle),
    .ap_ready(FloatvMultConst_15__ap_ready),
    .M(FloatvMultConst_15___M__q0),
    .P_N(FloatvMultConst_15___P_N__q0),
    .alpha_u(FloatvMultConst_15___alpha_u__q0),
    .fifo_in_s_dout(fifo_C_ch_result_Sextans_7__dout),
    .fifo_in_peek_dout(fifo_C_ch_result_Sextans_7__dout),
    .fifo_in_s_empty_n(fifo_C_ch_result_Sextans_7__empty_n),
    .fifo_in_peek_empty_n(fifo_C_ch_result_Sextans_7__empty_n),
    .fifo_in_s_read(fifo_C_ch_result_Sextans_7__read),
    .fifo_in_peek_read(),
    .fifo_out_din(fifo_C_ch_result_alpha_Sextans_7__din),
    .fifo_out_full_n(fifo_C_ch_result_alpha_Sextans_7__full_n),
    .fifo_out_write(fifo_C_ch_result_alpha_Sextans_7__write)
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_0__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_0__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_0__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_0__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_0__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_0__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_0__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_0__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_1__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_1__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_1__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_1__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_1__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_1__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_1__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_1__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_2__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_2__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_2__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_2__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_2__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_3__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_3__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_3__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_3__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_3__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_2__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_2__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_2__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_2__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_4__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_4__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_4__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_4__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_4__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_5__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_5__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_5__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_5__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_5__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_3__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_3__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_3__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_3__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_6__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_6__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_6__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_6__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_6__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_7__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_7__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_7__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_7__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_7__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_4__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_4__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_4__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_4__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_8__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_8__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_8__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_8__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_8__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_9__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_9__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_9__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_9__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_9__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_5__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_5__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_5__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_5__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_10__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_10__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_10__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_10__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_10__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_11__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_11__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_11__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_11__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_11__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_6__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_6__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_6__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_6__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_12__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_12__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_12__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_12__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_12__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_13__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_13__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_13__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_13__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_13__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) Merger
  Merger_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Merger_7__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_out_din(fifo_C_ch_result_Sextans_7__din),
    .fifo_out_full_n(fifo_C_ch_result_Sextans_7__full_n),
    .fifo_out_write(fifo_C_ch_result_Sextans_7__write),
    .fifo_in_0_dout(fifo_C_pe_Sextans_14__dout),
    .fifo_in_peek_0_dout(fifo_C_pe_Sextans_14__dout),
    .fifo_in_0_empty_n(fifo_C_pe_Sextans_14__empty_n),
    .fifo_in_peek_0_empty_n(fifo_C_pe_Sextans_14__empty_n),
    .fifo_in_0_read(fifo_C_pe_Sextans_14__read),
    .fifo_in_peek_0_read(),
    .fifo_in_1_dout(fifo_C_pe_Sextans_15__dout),
    .fifo_in_peek_1_dout(fifo_C_pe_Sextans_15__dout),
    .fifo_in_1_empty_n(fifo_C_pe_Sextans_15__empty_n),
    .fifo_in_peek_1_empty_n(fifo_C_pe_Sextans_15__empty_n),
    .fifo_in_1_read(fifo_C_pe_Sextans_15__read),
    .fifo_in_peek_1_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_0__ap_start),
    .ap_done(PEG_Bmtx_0__ap_done),
    .ap_idle(PEG_Bmtx_0__ap_idle),
    .ap_ready(PEG_Bmtx_0__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_0__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_0__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_0__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_0__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_0__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_1__din),
    .PE_inst_out_full_n(PE_inst_Sextans_1__full_n),
    .PE_inst_out_write(PE_inst_Sextans_1__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_0__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_0__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_0__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_0__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_0__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_0__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_0__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_0__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_0__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_0__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_0__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_0__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_0__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_1__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_1__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_1__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_1__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_1__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_2__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_2__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_2__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_2__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_2__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_3__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_3__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_3__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_3__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_3__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_4__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_4__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_4__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_5__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_5__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_5__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_6__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_6__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_6__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_7__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_7__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_7__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_0__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_0__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_0__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_1__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_1__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_1__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_2__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_2__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_2__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_3__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_3__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_3__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_0__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_0__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_0__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_0__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_0__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_1__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_1__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_1__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_0__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_0__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_0__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_1__ap_start),
    .ap_done(PEG_Bmtx_1__ap_done),
    .ap_idle(PEG_Bmtx_1__ap_idle),
    .ap_ready(PEG_Bmtx_1__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_1__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_1__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_1__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_1__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_1__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_2__din),
    .PE_inst_out_full_n(PE_inst_Sextans_2__full_n),
    .PE_inst_out_write(PE_inst_Sextans_2__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_1__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_1__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_1__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_1__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_1__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_1__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_1__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_1__read),
    .fifo_A_peek_read(),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_10__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_10__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_10__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_11__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_11__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_11__write),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_4__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_4__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_4__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_4__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_4__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_5__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_5__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_5__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_5__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_5__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_6__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_6__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_6__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_6__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_6__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_7__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_7__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_7__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_7__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_7__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_8__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_8__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_8__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_9__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_9__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_9__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_4__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_4__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_4__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_5__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_5__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_5__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_6__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_6__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_6__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_7__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_7__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_7__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_1__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_1__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_1__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_1__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_1__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_2__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_2__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_2__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_1__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_1__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_1__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_2__ap_start),
    .ap_done(PEG_Bmtx_2__ap_done),
    .ap_idle(PEG_Bmtx_2__ap_idle),
    .ap_ready(PEG_Bmtx_2__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_2__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_2__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_2__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_2__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_2__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_3__din),
    .PE_inst_out_full_n(PE_inst_Sextans_3__full_n),
    .PE_inst_out_write(PE_inst_Sextans_3__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_2__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_2__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_2__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_2__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_2__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_2__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_2__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_2__read),
    .fifo_A_peek_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_10__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_10__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_10__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_10__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_10__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_11__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_11__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_11__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_11__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_11__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_12__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_12__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_12__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_13__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_13__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_13__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_14__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_14__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_14__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_15__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_15__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_15__write),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_8__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_8__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_8__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_8__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_8__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_9__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_9__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_9__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_9__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_9__read),
    .fifo_B_in_peek_1_read(),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_10__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_10__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_10__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_11__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_11__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_11__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_8__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_8__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_8__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_9__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_9__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_9__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_2__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_2__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_2__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_2__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_2__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_3__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_3__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_3__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_2__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_2__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_2__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_3__ap_start),
    .ap_done(PEG_Bmtx_3__ap_done),
    .ap_idle(PEG_Bmtx_3__ap_idle),
    .ap_ready(PEG_Bmtx_3__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_3__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_3__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_3__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_3__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_3__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_4__din),
    .PE_inst_out_full_n(PE_inst_Sextans_4__full_n),
    .PE_inst_out_write(PE_inst_Sextans_4__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_3__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_3__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_3__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_3__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_3__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_3__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_3__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_3__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_12__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_12__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_12__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_12__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_12__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_13__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_13__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_13__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_13__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_13__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_14__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_14__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_14__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_14__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_14__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_15__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_15__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_15__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_15__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_15__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_16__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_16__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_16__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_17__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_17__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_17__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_18__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_18__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_18__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_19__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_19__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_19__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_12__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_12__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_12__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_13__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_13__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_13__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_14__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_14__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_14__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_15__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_15__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_15__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_3__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_3__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_3__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_3__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_3__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_4__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_4__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_4__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_3__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_3__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_3__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_4__ap_start),
    .ap_done(PEG_Bmtx_4__ap_done),
    .ap_idle(PEG_Bmtx_4__ap_idle),
    .ap_ready(PEG_Bmtx_4__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_4__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_4__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_4__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_4__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_4__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_5__din),
    .PE_inst_out_full_n(PE_inst_Sextans_5__full_n),
    .PE_inst_out_write(PE_inst_Sextans_5__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_4__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_4__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_4__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_4__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_4__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_4__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_4__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_4__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_16__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_16__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_16__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_16__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_16__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_17__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_17__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_17__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_17__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_17__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_18__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_18__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_18__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_18__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_18__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_19__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_19__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_19__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_19__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_19__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_20__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_20__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_20__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_21__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_21__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_21__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_22__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_22__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_22__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_23__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_23__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_23__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_16__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_16__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_16__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_17__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_17__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_17__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_18__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_18__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_18__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_19__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_19__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_19__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_4__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_4__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_4__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_4__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_4__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_5__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_5__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_5__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_4__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_4__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_4__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_5__ap_start),
    .ap_done(PEG_Bmtx_5__ap_done),
    .ap_idle(PEG_Bmtx_5__ap_idle),
    .ap_ready(PEG_Bmtx_5__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_5__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_5__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_5__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_5__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_5__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_6__din),
    .PE_inst_out_full_n(PE_inst_Sextans_6__full_n),
    .PE_inst_out_write(PE_inst_Sextans_6__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_5__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_5__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_5__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_5__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_5__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_5__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_5__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_5__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_20__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_20__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_20__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_20__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_20__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_21__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_21__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_21__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_21__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_21__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_22__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_22__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_22__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_22__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_22__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_23__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_23__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_23__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_23__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_23__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_24__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_24__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_24__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_25__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_25__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_25__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_26__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_26__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_26__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_27__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_27__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_27__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_20__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_20__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_20__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_21__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_21__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_21__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_22__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_22__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_22__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_23__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_23__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_23__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_5__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_5__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_5__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_5__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_5__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_6__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_6__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_6__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_5__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_5__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_5__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_6__ap_start),
    .ap_done(PEG_Bmtx_6__ap_done),
    .ap_idle(PEG_Bmtx_6__ap_idle),
    .ap_ready(PEG_Bmtx_6__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_6__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_6__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_6__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_6__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_6__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_7__din),
    .PE_inst_out_full_n(PE_inst_Sextans_7__full_n),
    .PE_inst_out_write(PE_inst_Sextans_7__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_6__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_6__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_6__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_6__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_6__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_6__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_6__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_6__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_24__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_24__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_24__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_24__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_24__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_25__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_25__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_25__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_25__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_25__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_26__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_26__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_26__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_26__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_26__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_27__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_27__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_27__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_27__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_27__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_28__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_28__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_28__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_29__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_29__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_29__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_30__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_30__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_30__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_31__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_31__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_31__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_24__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_24__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_24__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_25__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_25__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_25__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_26__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_26__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_26__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_27__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_27__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_27__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_6__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_6__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_6__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_6__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_6__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_7__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_7__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_7__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_6__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_6__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_6__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_7__ap_start),
    .ap_done(PEG_Bmtx_7__ap_done),
    .ap_idle(PEG_Bmtx_7__ap_idle),
    .ap_ready(PEG_Bmtx_7__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_7__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_7__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_7__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_7__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_7__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_8__din),
    .PE_inst_out_full_n(PE_inst_Sextans_8__full_n),
    .PE_inst_out_write(PE_inst_Sextans_8__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_7__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_7__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_7__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_7__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_7__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_7__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_7__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_7__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_28__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_28__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_28__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_28__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_28__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_29__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_29__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_29__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_29__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_29__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_30__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_30__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_30__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_30__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_30__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_31__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_31__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_31__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_31__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_31__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_32__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_32__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_32__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_33__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_33__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_33__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_34__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_34__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_34__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_35__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_35__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_35__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_28__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_28__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_28__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_29__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_29__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_29__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_30__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_30__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_30__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_31__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_31__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_31__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_7__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_7__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_7__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_7__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_7__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_8__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_8__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_8__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_7__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_7__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_7__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_8__ap_start),
    .ap_done(PEG_Bmtx_8__ap_done),
    .ap_idle(PEG_Bmtx_8__ap_idle),
    .ap_ready(PEG_Bmtx_8__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_8__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_8__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_8__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_8__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_8__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_9__din),
    .PE_inst_out_full_n(PE_inst_Sextans_9__full_n),
    .PE_inst_out_write(PE_inst_Sextans_9__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_8__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_8__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_8__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_8__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_8__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_8__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_8__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_8__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_32__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_32__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_32__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_32__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_32__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_33__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_33__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_33__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_33__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_33__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_34__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_34__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_34__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_34__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_34__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_35__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_35__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_35__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_35__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_35__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_36__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_36__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_36__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_37__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_37__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_37__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_38__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_38__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_38__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_39__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_39__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_39__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_32__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_32__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_32__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_33__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_33__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_33__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_34__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_34__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_34__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_35__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_35__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_35__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_8__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_8__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_8__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_8__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_8__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_9__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_9__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_9__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_8__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_8__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_8__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_9__ap_start),
    .ap_done(PEG_Bmtx_9__ap_done),
    .ap_idle(PEG_Bmtx_9__ap_idle),
    .ap_ready(PEG_Bmtx_9__ap_ready),
    .PE_inst_out_din(PE_inst_Sextans_10__din),
    .PE_inst_out_full_n(PE_inst_Sextans_10__full_n),
    .PE_inst_out_write(PE_inst_Sextans_10__write),
    .PE_inst_in_s_dout(PE_inst_Sextans_9__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_9__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_9__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_9__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_9__read),
    .PE_inst_in_peek_read(),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_9__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_9__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_9__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_9__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_9__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_9__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_9__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_9__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_36__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_36__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_36__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_36__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_36__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_37__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_37__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_37__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_37__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_37__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_38__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_38__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_38__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_38__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_38__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_39__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_39__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_39__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_39__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_39__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_40__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_40__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_40__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_41__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_41__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_41__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_42__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_42__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_42__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_43__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_43__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_43__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_36__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_36__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_36__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_37__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_37__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_37__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_38__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_38__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_38__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_39__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_39__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_39__write),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_10__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_10__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_10__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_9__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_9__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_9__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_9__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_9__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_9__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_9__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_9__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_10__ap_start),
    .ap_done(PEG_Bmtx_10__ap_done),
    .ap_idle(PEG_Bmtx_10__ap_idle),
    .ap_ready(PEG_Bmtx_10__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_10__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_10__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_10__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_10__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_10__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_11__din),
    .PE_inst_out_full_n(PE_inst_Sextans_11__full_n),
    .PE_inst_out_write(PE_inst_Sextans_11__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_10__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_10__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_10__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_10__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_10__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_10__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_10__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_10__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_40__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_40__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_40__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_40__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_40__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_41__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_41__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_41__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_41__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_41__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_42__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_42__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_42__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_42__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_42__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_43__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_43__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_43__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_43__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_43__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_44__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_44__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_44__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_45__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_45__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_45__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_46__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_46__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_46__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_47__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_47__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_47__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_40__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_40__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_40__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_41__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_41__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_41__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_42__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_42__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_42__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_43__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_43__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_43__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_10__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_10__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_10__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_10__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_10__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_11__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_11__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_11__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_10__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_10__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_10__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_11__ap_start),
    .ap_done(PEG_Bmtx_11__ap_done),
    .ap_idle(PEG_Bmtx_11__ap_idle),
    .ap_ready(PEG_Bmtx_11__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_11__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_11__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_11__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_11__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_11__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_12__din),
    .PE_inst_out_full_n(PE_inst_Sextans_12__full_n),
    .PE_inst_out_write(PE_inst_Sextans_12__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_11__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_11__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_11__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_11__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_11__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_11__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_11__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_11__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_44__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_44__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_44__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_44__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_44__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_45__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_45__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_45__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_45__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_45__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_46__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_46__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_46__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_46__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_46__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_47__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_47__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_47__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_47__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_47__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_48__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_48__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_48__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_49__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_49__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_49__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_50__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_50__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_50__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_51__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_51__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_51__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_44__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_44__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_44__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_45__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_45__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_45__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_46__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_46__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_46__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_47__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_47__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_47__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_11__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_11__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_11__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_11__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_11__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_12__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_12__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_12__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_11__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_11__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_11__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_12__ap_start),
    .ap_done(PEG_Bmtx_12__ap_done),
    .ap_idle(PEG_Bmtx_12__ap_idle),
    .ap_ready(PEG_Bmtx_12__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_12__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_12__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_12__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_12__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_12__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_13__din),
    .PE_inst_out_full_n(PE_inst_Sextans_13__full_n),
    .PE_inst_out_write(PE_inst_Sextans_13__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_12__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_12__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_12__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_12__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_12__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_12__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_12__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_12__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_48__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_48__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_48__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_48__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_48__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_49__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_49__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_49__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_49__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_49__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_50__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_50__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_50__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_50__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_50__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_51__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_51__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_51__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_51__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_51__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_52__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_52__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_52__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_53__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_53__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_53__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_54__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_54__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_54__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_55__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_55__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_55__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_48__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_48__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_48__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_49__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_49__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_49__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_50__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_50__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_50__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_51__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_51__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_51__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_12__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_12__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_12__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_12__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_12__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_13__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_13__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_13__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_12__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_12__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_12__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_13__ap_start),
    .ap_done(PEG_Bmtx_13__ap_done),
    .ap_idle(PEG_Bmtx_13__ap_idle),
    .ap_ready(PEG_Bmtx_13__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_13__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_13__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_13__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_13__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_13__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_14__din),
    .PE_inst_out_full_n(PE_inst_Sextans_14__full_n),
    .PE_inst_out_write(PE_inst_Sextans_14__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_13__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_13__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_13__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_13__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_13__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_13__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_13__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_13__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_52__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_52__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_52__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_52__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_52__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_53__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_53__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_53__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_53__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_53__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_54__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_54__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_54__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_54__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_54__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_55__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_55__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_55__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_55__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_55__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_56__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_56__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_56__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_57__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_57__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_57__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_58__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_58__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_58__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_59__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_59__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_59__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_52__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_52__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_52__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_53__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_53__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_53__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_54__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_54__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_54__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_55__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_55__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_55__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_13__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_13__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_13__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_13__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_13__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_14__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_14__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_14__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_13__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_13__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_13__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_14__ap_start),
    .ap_done(PEG_Bmtx_14__ap_done),
    .ap_idle(PEG_Bmtx_14__ap_idle),
    .ap_ready(PEG_Bmtx_14__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_14__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_14__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_14__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_14__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_14__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_15__din),
    .PE_inst_out_full_n(PE_inst_Sextans_15__full_n),
    .PE_inst_out_write(PE_inst_Sextans_15__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_14__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_14__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_14__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_14__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_14__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_14__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_14__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_14__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_56__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_56__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_56__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_56__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_56__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_57__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_57__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_57__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_57__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_57__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_58__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_58__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_58__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_58__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_58__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_59__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_59__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_59__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_59__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_59__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_60__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_60__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_60__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_61__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_61__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_61__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_62__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_62__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_62__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_63__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_63__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_63__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_56__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_56__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_56__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_57__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_57__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_57__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_58__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_58__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_58__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_59__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_59__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_59__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_14__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_14__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_14__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_14__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_14__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_15__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_15__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_15__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_14__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_14__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_14__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Bmtx
  PEG_Bmtx_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Bmtx_15__ap_start),
    .ap_done(PEG_Bmtx_15__ap_done),
    .ap_idle(PEG_Bmtx_15__ap_idle),
    .ap_ready(PEG_Bmtx_15__ap_ready),
    .PE_inst_in_s_dout(PE_inst_Sextans_15__dout),
    .PE_inst_in_peek_dout(PE_inst_Sextans_15__dout),
    .PE_inst_in_s_empty_n(PE_inst_Sextans_15__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_Sextans_15__empty_n),
    .PE_inst_in_s_read(PE_inst_Sextans_15__read),
    .PE_inst_in_peek_read(),
    .PE_inst_out_din(PE_inst_Sextans_16__din),
    .PE_inst_out_full_n(PE_inst_Sextans_16__full_n),
    .PE_inst_out_write(PE_inst_Sextans_16__write),
    .PE_inst_to_Cmtx_din(PE_inst_to_Cmtx_Sextans_15__din),
    .PE_inst_to_Cmtx_full_n(PE_inst_to_Cmtx_Sextans_15__full_n),
    .PE_inst_to_Cmtx_write(PE_inst_to_Cmtx_Sextans_15__write),
    .fifo_A_s_dout(fifo_A_pe_Sextans_15__dout),
    .fifo_A_peek_dout(fifo_A_pe_Sextans_15__dout),
    .fifo_A_s_empty_n(fifo_A_pe_Sextans_15__empty_n),
    .fifo_A_peek_empty_n(fifo_A_pe_Sextans_15__empty_n),
    .fifo_A_s_read(fifo_A_pe_Sextans_15__read),
    .fifo_A_peek_read(),
    .fifo_B_in_0_dout(fifo_B_pe_Sextans_60__dout),
    .fifo_B_in_peek_0_dout(fifo_B_pe_Sextans_60__dout),
    .fifo_B_in_0_empty_n(fifo_B_pe_Sextans_60__empty_n),
    .fifo_B_in_peek_0_empty_n(fifo_B_pe_Sextans_60__empty_n),
    .fifo_B_in_0_read(fifo_B_pe_Sextans_60__read),
    .fifo_B_in_peek_0_read(),
    .fifo_B_in_1_dout(fifo_B_pe_Sextans_61__dout),
    .fifo_B_in_peek_1_dout(fifo_B_pe_Sextans_61__dout),
    .fifo_B_in_1_empty_n(fifo_B_pe_Sextans_61__empty_n),
    .fifo_B_in_peek_1_empty_n(fifo_B_pe_Sextans_61__empty_n),
    .fifo_B_in_1_read(fifo_B_pe_Sextans_61__read),
    .fifo_B_in_peek_1_read(),
    .fifo_B_in_2_dout(fifo_B_pe_Sextans_62__dout),
    .fifo_B_in_peek_2_dout(fifo_B_pe_Sextans_62__dout),
    .fifo_B_in_2_empty_n(fifo_B_pe_Sextans_62__empty_n),
    .fifo_B_in_peek_2_empty_n(fifo_B_pe_Sextans_62__empty_n),
    .fifo_B_in_2_read(fifo_B_pe_Sextans_62__read),
    .fifo_B_in_peek_2_read(),
    .fifo_B_in_3_dout(fifo_B_pe_Sextans_63__dout),
    .fifo_B_in_peek_3_dout(fifo_B_pe_Sextans_63__dout),
    .fifo_B_in_3_empty_n(fifo_B_pe_Sextans_63__empty_n),
    .fifo_B_in_peek_3_empty_n(fifo_B_pe_Sextans_63__empty_n),
    .fifo_B_in_3_read(fifo_B_pe_Sextans_63__read),
    .fifo_B_in_peek_3_read(),
    .fifo_B_out_0_din(fifo_B_pe_Sextans_64__din),
    .fifo_B_out_0_full_n(fifo_B_pe_Sextans_64__full_n),
    .fifo_B_out_0_write(fifo_B_pe_Sextans_64__write),
    .fifo_B_out_1_din(fifo_B_pe_Sextans_65__din),
    .fifo_B_out_1_full_n(fifo_B_pe_Sextans_65__full_n),
    .fifo_B_out_1_write(fifo_B_pe_Sextans_65__write),
    .fifo_B_out_2_din(fifo_B_pe_Sextans_66__din),
    .fifo_B_out_2_full_n(fifo_B_pe_Sextans_66__full_n),
    .fifo_B_out_2_write(fifo_B_pe_Sextans_66__write),
    .fifo_B_out_3_din(fifo_B_pe_Sextans_67__din),
    .fifo_B_out_3_full_n(fifo_B_pe_Sextans_67__full_n),
    .fifo_B_out_3_write(fifo_B_pe_Sextans_67__write),
    .fifo_aBvec_0_din(fifo_aBvec_Sextans_60__din),
    .fifo_aBvec_0_full_n(fifo_aBvec_Sextans_60__full_n),
    .fifo_aBvec_0_write(fifo_aBvec_Sextans_60__write),
    .fifo_aBvec_1_din(fifo_aBvec_Sextans_61__din),
    .fifo_aBvec_1_full_n(fifo_aBvec_Sextans_61__full_n),
    .fifo_aBvec_1_write(fifo_aBvec_Sextans_61__write),
    .fifo_aBvec_2_din(fifo_aBvec_Sextans_62__din),
    .fifo_aBvec_2_full_n(fifo_aBvec_Sextans_62__full_n),
    .fifo_aBvec_2_write(fifo_aBvec_Sextans_62__write),
    .fifo_aBvec_3_din(fifo_aBvec_Sextans_63__din),
    .fifo_aBvec_3_full_n(fifo_aBvec_Sextans_63__full_n),
    .fifo_aBvec_3_write(fifo_aBvec_Sextans_63__write),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_Sextans_15__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_Sextans_15__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_Sextans_15__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_Sextans_15__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_Sextans_15__read),
    .fifo_inst_in_peek_read(),
    .fifo_inst_out_din(fifo_edge_list_ptr_Sextans_16__din),
    .fifo_inst_out_full_n(fifo_edge_list_ptr_Sextans_16__full_n),
    .fifo_inst_out_write(fifo_edge_list_ptr_Sextans_16__write),
    .fifo_inst_out_to_Cmtx_din(fifo_edge_list_ptr_to_Cmtx_Sextans_15__din),
    .fifo_inst_out_to_Cmtx_full_n(fifo_edge_list_ptr_to_Cmtx_Sextans_15__full_n),
    .fifo_inst_out_to_Cmtx_write(fifo_edge_list_ptr_to_Cmtx_Sextans_15__write)
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_0__ap_start),
    .ap_done(PEG_Cmtx_0__ap_done),
    .ap_idle(PEG_Cmtx_0__ap_idle),
    .ap_ready(PEG_Cmtx_0__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_0__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_0__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_0__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_0__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_0__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_0__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_0__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_0__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_0__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_0__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_0__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_0__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_0__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_1__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_1__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_1__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_1__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_1__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_2__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_2__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_2__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_2__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_2__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_3__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_3__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_3__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_3__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_3__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_0__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_0__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_0__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_0__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_0__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_1__ap_start),
    .ap_done(PEG_Cmtx_1__ap_done),
    .ap_idle(PEG_Cmtx_1__ap_idle),
    .ap_ready(PEG_Cmtx_1__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_1__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_1__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_1__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_1__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_1__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_1__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_1__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_1__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_4__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_4__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_4__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_4__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_4__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_5__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_5__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_5__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_5__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_5__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_6__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_6__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_6__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_6__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_6__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_7__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_7__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_7__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_7__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_7__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_1__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_1__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_1__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_1__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_1__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_2__ap_start),
    .ap_done(PEG_Cmtx_2__ap_done),
    .ap_idle(PEG_Cmtx_2__ap_idle),
    .ap_ready(PEG_Cmtx_2__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_2__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_2__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_2__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_2__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_2__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_2__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_2__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_2__write),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_10__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_10__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_10__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_10__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_10__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_11__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_11__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_11__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_11__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_11__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_8__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_8__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_8__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_8__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_8__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_9__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_9__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_9__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_9__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_9__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_2__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_2__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_2__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_2__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_2__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_3__ap_start),
    .ap_done(PEG_Cmtx_3__ap_done),
    .ap_idle(PEG_Cmtx_3__ap_idle),
    .ap_ready(PEG_Cmtx_3__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_3__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_3__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_3__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_3__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_3__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_3__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_3__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_3__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_12__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_12__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_12__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_12__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_12__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_13__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_13__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_13__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_13__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_13__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_14__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_14__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_14__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_14__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_14__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_15__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_15__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_15__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_15__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_15__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_3__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_3__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_3__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_3__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_3__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_4__ap_start),
    .ap_done(PEG_Cmtx_4__ap_done),
    .ap_idle(PEG_Cmtx_4__ap_idle),
    .ap_ready(PEG_Cmtx_4__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_4__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_4__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_4__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_4__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_4__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_4__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_4__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_4__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_16__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_16__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_16__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_16__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_16__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_17__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_17__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_17__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_17__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_17__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_18__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_18__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_18__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_18__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_18__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_19__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_19__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_19__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_19__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_19__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_4__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_4__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_4__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_4__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_4__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_5__ap_start),
    .ap_done(PEG_Cmtx_5__ap_done),
    .ap_idle(PEG_Cmtx_5__ap_idle),
    .ap_ready(PEG_Cmtx_5__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_5__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_5__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_5__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_5__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_5__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_5__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_5__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_5__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_20__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_20__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_20__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_20__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_20__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_21__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_21__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_21__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_21__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_21__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_22__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_22__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_22__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_22__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_22__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_23__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_23__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_23__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_23__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_23__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_5__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_5__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_5__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_5__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_5__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_6__ap_start),
    .ap_done(PEG_Cmtx_6__ap_done),
    .ap_idle(PEG_Cmtx_6__ap_idle),
    .ap_ready(PEG_Cmtx_6__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_6__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_6__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_6__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_6__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_6__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_6__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_6__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_6__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_24__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_24__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_24__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_24__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_24__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_25__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_25__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_25__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_25__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_25__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_26__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_26__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_26__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_26__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_26__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_27__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_27__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_27__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_27__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_27__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_6__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_6__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_6__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_6__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_6__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_7__ap_start),
    .ap_done(PEG_Cmtx_7__ap_done),
    .ap_idle(PEG_Cmtx_7__ap_idle),
    .ap_ready(PEG_Cmtx_7__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_7__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_7__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_7__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_7__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_7__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_7__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_7__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_7__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_28__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_28__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_28__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_28__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_28__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_29__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_29__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_29__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_29__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_29__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_30__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_30__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_30__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_30__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_30__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_31__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_31__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_31__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_31__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_31__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_7__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_7__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_7__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_7__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_7__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_8__ap_start),
    .ap_done(PEG_Cmtx_8__ap_done),
    .ap_idle(PEG_Cmtx_8__ap_idle),
    .ap_ready(PEG_Cmtx_8__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_8__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_8__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_8__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_8__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_8__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_8__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_8__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_8__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_32__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_32__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_32__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_32__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_32__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_33__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_33__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_33__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_33__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_33__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_34__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_34__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_34__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_34__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_34__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_35__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_35__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_35__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_35__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_35__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_8__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_8__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_8__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_8__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_8__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_9__ap_start),
    .ap_done(PEG_Cmtx_9__ap_done),
    .ap_idle(PEG_Cmtx_9__ap_idle),
    .ap_ready(PEG_Cmtx_9__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_9__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_9__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_9__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_9__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_9__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_9__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_9__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_9__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_36__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_36__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_36__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_36__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_36__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_37__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_37__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_37__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_37__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_37__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_38__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_38__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_38__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_38__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_38__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_39__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_39__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_39__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_39__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_39__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_9__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_9__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_9__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_9__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_9__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_10__ap_start),
    .ap_done(PEG_Cmtx_10__ap_done),
    .ap_idle(PEG_Cmtx_10__ap_idle),
    .ap_ready(PEG_Cmtx_10__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_10__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_10__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_10__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_10__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_10__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_10__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_10__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_10__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_40__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_40__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_40__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_40__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_40__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_41__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_41__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_41__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_41__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_41__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_42__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_42__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_42__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_42__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_42__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_43__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_43__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_43__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_43__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_43__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_10__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_10__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_10__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_10__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_10__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_11__ap_start),
    .ap_done(PEG_Cmtx_11__ap_done),
    .ap_idle(PEG_Cmtx_11__ap_idle),
    .ap_ready(PEG_Cmtx_11__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_11__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_11__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_11__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_11__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_11__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_11__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_11__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_11__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_44__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_44__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_44__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_44__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_44__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_45__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_45__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_45__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_45__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_45__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_46__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_46__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_46__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_46__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_46__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_47__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_47__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_47__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_47__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_47__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_11__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_11__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_11__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_11__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_11__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_12__ap_start),
    .ap_done(PEG_Cmtx_12__ap_done),
    .ap_idle(PEG_Cmtx_12__ap_idle),
    .ap_ready(PEG_Cmtx_12__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_12__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_12__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_12__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_12__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_12__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_12__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_12__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_12__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_48__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_48__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_48__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_48__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_48__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_49__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_49__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_49__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_49__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_49__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_50__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_50__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_50__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_50__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_50__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_51__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_51__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_51__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_51__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_51__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_12__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_12__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_12__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_12__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_12__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_13__ap_start),
    .ap_done(PEG_Cmtx_13__ap_done),
    .ap_idle(PEG_Cmtx_13__ap_idle),
    .ap_ready(PEG_Cmtx_13__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_13__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_13__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_13__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_13__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_13__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_13__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_13__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_13__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_52__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_52__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_52__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_52__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_52__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_53__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_53__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_53__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_53__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_53__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_54__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_54__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_54__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_54__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_54__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_55__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_55__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_55__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_55__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_55__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_13__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_13__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_13__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_13__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_13__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_14__ap_start),
    .ap_done(PEG_Cmtx_14__ap_done),
    .ap_idle(PEG_Cmtx_14__ap_idle),
    .ap_ready(PEG_Cmtx_14__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_14__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_14__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_14__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_14__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_14__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_14__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_14__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_14__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_56__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_56__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_56__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_56__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_56__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_57__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_57__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_57__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_57__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_57__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_58__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_58__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_58__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_58__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_58__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_59__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_59__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_59__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_59__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_59__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_14__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_14__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_14__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_14__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_14__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PEG_Cmtx
  PEG_Cmtx_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PEG_Cmtx_15__ap_start),
    .ap_done(PEG_Cmtx_15__ap_done),
    .ap_idle(PEG_Cmtx_15__ap_idle),
    .ap_ready(PEG_Cmtx_15__ap_ready),
    .PE_inst_in_s_dout(PE_inst_to_Cmtx_Sextans_15__dout),
    .PE_inst_in_peek_dout(PE_inst_to_Cmtx_Sextans_15__dout),
    .PE_inst_in_s_empty_n(PE_inst_to_Cmtx_Sextans_15__empty_n),
    .PE_inst_in_peek_empty_n(PE_inst_to_Cmtx_Sextans_15__empty_n),
    .PE_inst_in_s_read(PE_inst_to_Cmtx_Sextans_15__read),
    .PE_inst_in_peek_read(),
    .fifo_C_out_din(fifo_C_pe_Sextans_15__din),
    .fifo_C_out_full_n(fifo_C_pe_Sextans_15__full_n),
    .fifo_C_out_write(fifo_C_pe_Sextans_15__write),
    .fifo_aBvec_0_dout(fifo_aBvec_Sextans_60__dout),
    .fifo_aBvec_peek_0_dout(fifo_aBvec_Sextans_60__dout),
    .fifo_aBvec_0_empty_n(fifo_aBvec_Sextans_60__empty_n),
    .fifo_aBvec_peek_0_empty_n(fifo_aBvec_Sextans_60__empty_n),
    .fifo_aBvec_0_read(fifo_aBvec_Sextans_60__read),
    .fifo_aBvec_peek_0_read(),
    .fifo_aBvec_1_dout(fifo_aBvec_Sextans_61__dout),
    .fifo_aBvec_peek_1_dout(fifo_aBvec_Sextans_61__dout),
    .fifo_aBvec_1_empty_n(fifo_aBvec_Sextans_61__empty_n),
    .fifo_aBvec_peek_1_empty_n(fifo_aBvec_Sextans_61__empty_n),
    .fifo_aBvec_1_read(fifo_aBvec_Sextans_61__read),
    .fifo_aBvec_peek_1_read(),
    .fifo_aBvec_2_dout(fifo_aBvec_Sextans_62__dout),
    .fifo_aBvec_peek_2_dout(fifo_aBvec_Sextans_62__dout),
    .fifo_aBvec_2_empty_n(fifo_aBvec_Sextans_62__empty_n),
    .fifo_aBvec_peek_2_empty_n(fifo_aBvec_Sextans_62__empty_n),
    .fifo_aBvec_2_read(fifo_aBvec_Sextans_62__read),
    .fifo_aBvec_peek_2_read(),
    .fifo_aBvec_3_dout(fifo_aBvec_Sextans_63__dout),
    .fifo_aBvec_peek_3_dout(fifo_aBvec_Sextans_63__dout),
    .fifo_aBvec_3_empty_n(fifo_aBvec_Sextans_63__empty_n),
    .fifo_aBvec_peek_3_empty_n(fifo_aBvec_Sextans_63__empty_n),
    .fifo_aBvec_3_read(fifo_aBvec_Sextans_63__read),
    .fifo_aBvec_peek_3_read(),
    .fifo_inst_in_s_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_15__dout),
    .fifo_inst_in_peek_dout(fifo_edge_list_ptr_to_Cmtx_Sextans_15__dout),
    .fifo_inst_in_s_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_15__empty_n),
    .fifo_inst_in_peek_empty_n(fifo_edge_list_ptr_to_Cmtx_Sextans_15__empty_n),
    .fifo_inst_in_s_read(fifo_edge_list_ptr_to_Cmtx_Sextans_15__read),
    .fifo_inst_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_0__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_0__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_0__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_0__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_0__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_0__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_0__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_0__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_1__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_1__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_1__write)
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_1__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_1__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_1__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_1__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_1__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_2__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_2__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_2__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_3__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_3__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_3__write)
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_2__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_2__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_2__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_2__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_2__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_2__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_4__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_4__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_4__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_5__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_5__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_5__write)
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_3__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_3__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_3__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_3__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_3__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_3__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_6__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_6__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_6__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_7__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_7__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_7__write)
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_4__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_4__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_4__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_4__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_4__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_4__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_8__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_8__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_8__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_9__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_9__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_9__write)
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_5__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_5__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_5__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_5__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_5__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_5__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_10__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_10__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_10__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_11__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_11__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_11__write)
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_6__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_6__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_6__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_6__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_6__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_6__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_12__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_12__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_12__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_13__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_13__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_13__write)
  );


  (* keep_hierarchy = "yes" *) Scatter_1_2
  Scatter_1_2_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Scatter_1_2_7__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_A_Sextans_7__dout),
    .fifo_in_peek_dout(fifo_A_Sextans_7__dout),
    .fifo_in_s_empty_n(fifo_A_Sextans_7__empty_n),
    .fifo_in_peek_empty_n(fifo_A_Sextans_7__empty_n),
    .fifo_in_s_read(fifo_A_Sextans_7__read),
    .fifo_in_peek_read(),
    .fifo_out_0_din(fifo_A_pe_Sextans_14__din),
    .fifo_out_0_full_n(fifo_A_pe_Sextans_14__full_n),
    .fifo_out_0_write(fifo_A_pe_Sextans_14__write),
    .fifo_out_1_din(fifo_A_pe_Sextans_15__din),
    .fifo_out_1_full_n(fifo_A_pe_Sextans_15__full_n),
    .fifo_out_1_write(fifo_A_pe_Sextans_15__write)
  );


  (* keep_hierarchy = "yes" *) black_hole_float_v16
  black_hole_float_v16_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(black_hole_float_v16_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_B_pe_Sextans_64__dout),
    .fifo_in_peek_dout(fifo_B_pe_Sextans_64__dout),
    .fifo_in_s_empty_n(fifo_B_pe_Sextans_64__empty_n),
    .fifo_in_peek_empty_n(fifo_B_pe_Sextans_64__empty_n),
    .fifo_in_s_read(fifo_B_pe_Sextans_64__read),
    .fifo_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) black_hole_float_v16
  black_hole_float_v16_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(black_hole_float_v16_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_B_pe_Sextans_65__dout),
    .fifo_in_peek_dout(fifo_B_pe_Sextans_65__dout),
    .fifo_in_s_empty_n(fifo_B_pe_Sextans_65__empty_n),
    .fifo_in_peek_empty_n(fifo_B_pe_Sextans_65__empty_n),
    .fifo_in_s_read(fifo_B_pe_Sextans_65__read),
    .fifo_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) black_hole_float_v16
  black_hole_float_v16_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(black_hole_float_v16_2__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_B_pe_Sextans_66__dout),
    .fifo_in_peek_dout(fifo_B_pe_Sextans_66__dout),
    .fifo_in_s_empty_n(fifo_B_pe_Sextans_66__empty_n),
    .fifo_in_peek_empty_n(fifo_B_pe_Sextans_66__empty_n),
    .fifo_in_s_read(fifo_B_pe_Sextans_66__read),
    .fifo_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) black_hole_float_v16
  black_hole_float_v16_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(black_hole_float_v16_3__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_B_pe_Sextans_67__dout),
    .fifo_in_peek_dout(fifo_B_pe_Sextans_67__dout),
    .fifo_in_s_empty_n(fifo_B_pe_Sextans_67__empty_n),
    .fifo_in_peek_empty_n(fifo_B_pe_Sextans_67__empty_n),
    .fifo_in_s_read(fifo_B_pe_Sextans_67__read),
    .fifo_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) black_hole_int
  black_hole_int_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(black_hole_int_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(PE_inst_Sextans_16__dout),
    .fifo_in_peek_dout(PE_inst_Sextans_16__dout),
    .fifo_in_s_empty_n(PE_inst_Sextans_16__empty_n),
    .fifo_in_peek_empty_n(PE_inst_Sextans_16__empty_n),
    .fifo_in_s_read(PE_inst_Sextans_16__read),
    .fifo_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) black_hole_int
  black_hole_int_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(black_hole_int_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_in_s_dout(fifo_edge_list_ptr_Sextans_16__dout),
    .fifo_in_peek_dout(fifo_edge_list_ptr_Sextans_16__dout),
    .fifo_in_s_empty_n(fifo_edge_list_ptr_Sextans_16__empty_n),
    .fifo_in_peek_empty_n(fifo_edge_list_ptr_Sextans_16__empty_n),
    .fifo_in_s_read(fifo_edge_list_ptr_Sextans_16__read),
    .fifo_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_0__ap_start),
    .ap_done(read_A_0__ap_done),
    .ap_idle(read_A_0__ap_idle),
    .ap_ready(read_A_0__ap_ready),
    .A_len(read_A_0___NUM_A_LEN__q0),
    .P_N(read_A_0___P_N__q0),
    .A_read_addr_din(edge_list_ch_0_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_0_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_0_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_0_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_0_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_0_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_0_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_0_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_0_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_0_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_0_write_addr__write),
    .A_write_data_din(edge_list_ch_0_write_data__din),
    .A_write_data_full_n(edge_list_ch_0_write_data__full_n),
    .A_write_data_write(edge_list_ch_0_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_0_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_0_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_0_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_0_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_0_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_0__din),
    .fifo_A_full_n(fifo_A_Sextans_0__full_n),
    .fifo_A_write(fifo_A_Sextans_0__write)
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_1__ap_start),
    .ap_done(read_A_1__ap_done),
    .ap_idle(read_A_1__ap_idle),
    .ap_ready(read_A_1__ap_ready),
    .A_len(read_A_1___NUM_A_LEN__q0),
    .P_N(read_A_1___P_N__q0),
    .A_read_addr_din(edge_list_ch_1_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_1_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_1_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_1_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_1_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_1_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_1_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_1_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_1_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_1_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_1_write_addr__write),
    .A_write_data_din(edge_list_ch_1_write_data__din),
    .A_write_data_full_n(edge_list_ch_1_write_data__full_n),
    .A_write_data_write(edge_list_ch_1_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_1_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_1_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_1_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_1_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_1_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_1__din),
    .fifo_A_full_n(fifo_A_Sextans_1__full_n),
    .fifo_A_write(fifo_A_Sextans_1__write)
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_2__ap_start),
    .ap_done(read_A_2__ap_done),
    .ap_idle(read_A_2__ap_idle),
    .ap_ready(read_A_2__ap_ready),
    .A_len(read_A_2___NUM_A_LEN__q0),
    .P_N(read_A_2___P_N__q0),
    .A_read_addr_din(edge_list_ch_2_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_2_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_2_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_2_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_2_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_2_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_2_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_2_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_2_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_2_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_2_write_addr__write),
    .A_write_data_din(edge_list_ch_2_write_data__din),
    .A_write_data_full_n(edge_list_ch_2_write_data__full_n),
    .A_write_data_write(edge_list_ch_2_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_2_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_2_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_2_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_2_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_2_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_2__din),
    .fifo_A_full_n(fifo_A_Sextans_2__full_n),
    .fifo_A_write(fifo_A_Sextans_2__write)
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_3__ap_start),
    .ap_done(read_A_3__ap_done),
    .ap_idle(read_A_3__ap_idle),
    .ap_ready(read_A_3__ap_ready),
    .A_len(read_A_3___NUM_A_LEN__q0),
    .P_N(read_A_3___P_N__q0),
    .A_read_addr_din(edge_list_ch_3_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_3_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_3_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_3_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_3_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_3_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_3_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_3_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_3_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_3_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_3_write_addr__write),
    .A_write_data_din(edge_list_ch_3_write_data__din),
    .A_write_data_full_n(edge_list_ch_3_write_data__full_n),
    .A_write_data_write(edge_list_ch_3_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_3_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_3_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_3_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_3_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_3_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_3__din),
    .fifo_A_full_n(fifo_A_Sextans_3__full_n),
    .fifo_A_write(fifo_A_Sextans_3__write)
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_4__ap_start),
    .ap_done(read_A_4__ap_done),
    .ap_idle(read_A_4__ap_idle),
    .ap_ready(read_A_4__ap_ready),
    .A_len(read_A_4___NUM_A_LEN__q0),
    .P_N(read_A_4___P_N__q0),
    .A_read_addr_din(edge_list_ch_4_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_4_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_4_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_4_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_4_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_4_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_4_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_4_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_4_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_4_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_4_write_addr__write),
    .A_write_data_din(edge_list_ch_4_write_data__din),
    .A_write_data_full_n(edge_list_ch_4_write_data__full_n),
    .A_write_data_write(edge_list_ch_4_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_4_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_4_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_4_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_4_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_4_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_4__din),
    .fifo_A_full_n(fifo_A_Sextans_4__full_n),
    .fifo_A_write(fifo_A_Sextans_4__write)
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_5__ap_start),
    .ap_done(read_A_5__ap_done),
    .ap_idle(read_A_5__ap_idle),
    .ap_ready(read_A_5__ap_ready),
    .A_len(read_A_5___NUM_A_LEN__q0),
    .P_N(read_A_5___P_N__q0),
    .A_read_addr_din(edge_list_ch_5_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_5_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_5_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_5_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_5_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_5_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_5_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_5_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_5_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_5_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_5_write_addr__write),
    .A_write_data_din(edge_list_ch_5_write_data__din),
    .A_write_data_full_n(edge_list_ch_5_write_data__full_n),
    .A_write_data_write(edge_list_ch_5_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_5_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_5_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_5_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_5_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_5_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_5__din),
    .fifo_A_full_n(fifo_A_Sextans_5__full_n),
    .fifo_A_write(fifo_A_Sextans_5__write)
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_6__ap_start),
    .ap_done(read_A_6__ap_done),
    .ap_idle(read_A_6__ap_idle),
    .ap_ready(read_A_6__ap_ready),
    .A_len(read_A_6___NUM_A_LEN__q0),
    .P_N(read_A_6___P_N__q0),
    .A_read_addr_din(edge_list_ch_6_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_6_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_6_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_6_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_6_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_6_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_6_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_6_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_6_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_6_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_6_write_addr__write),
    .A_write_data_din(edge_list_ch_6_write_data__din),
    .A_write_data_full_n(edge_list_ch_6_write_data__full_n),
    .A_write_data_write(edge_list_ch_6_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_6_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_6_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_6_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_6_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_6_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_6__din),
    .fifo_A_full_n(fifo_A_Sextans_6__full_n),
    .fifo_A_write(fifo_A_Sextans_6__write)
  );


  (* keep_hierarchy = "yes" *) read_A
  read_A_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_A_7__ap_start),
    .ap_done(read_A_7__ap_done),
    .ap_idle(read_A_7__ap_idle),
    .ap_ready(read_A_7__ap_ready),
    .A_len(read_A_7___NUM_A_LEN__q0),
    .P_N(read_A_7___P_N__q0),
    .A_read_addr_din(edge_list_ch_7_read_addr__din),
    .A_read_addr_full_n(edge_list_ch_7_read_addr__full_n),
    .A_read_addr_write(edge_list_ch_7_read_addr__write),
    .A_read_data_s_dout({1'b0, edge_list_ch_7_read_data__dout}),
    .A_read_data_peek_dout({1'b0, edge_list_ch_7_read_data__dout}),
    .A_read_data_s_empty_n(edge_list_ch_7_read_data__empty_n),
    .A_read_data_peek_empty_n(edge_list_ch_7_read_data__empty_n),
    .A_read_data_s_read(edge_list_ch_7_read_data__read),
    .A_read_data_peek_read(),
    .A_write_addr_din(edge_list_ch_7_write_addr__din),
    .A_write_addr_full_n(edge_list_ch_7_write_addr__full_n),
    .A_write_addr_write(edge_list_ch_7_write_addr__write),
    .A_write_data_din(edge_list_ch_7_write_data__din),
    .A_write_data_full_n(edge_list_ch_7_write_data__full_n),
    .A_write_data_write(edge_list_ch_7_write_data__write),
    .A_write_resp_s_dout({1'b0, edge_list_ch_7_write_resp__dout}),
    .A_write_resp_peek_dout({1'b0, edge_list_ch_7_write_resp__dout}),
    .A_write_resp_s_empty_n(edge_list_ch_7_write_resp__empty_n),
    .A_write_resp_peek_empty_n(edge_list_ch_7_write_resp__empty_n),
    .A_write_resp_s_read(edge_list_ch_7_write_resp__read),
    .A_write_resp_peek_read(),
    .fifo_A_din(fifo_A_Sextans_7__din),
    .fifo_A_full_n(fifo_A_Sextans_7__full_n),
    .fifo_A_write(fifo_A_Sextans_7__write)
  );


  (* keep_hierarchy = "yes" *) read_B
  read_B_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_B_0__ap_start),
    .ap_done(read_B_0__ap_done),
    .ap_idle(read_B_0__ap_idle),
    .ap_ready(read_B_0__ap_ready),
    .K(read_B_0___K__q0),
    .P_N(read_B_0___P_N__q0),
    .fifo_B_din(fifo_B_pe_Sextans_0__din),
    .fifo_B_full_n(fifo_B_pe_Sextans_0__full_n),
    .fifo_B_write(fifo_B_pe_Sextans_0__write),
    .B_read_addr_din(mat_B_ch_0_read_addr__din),
    .B_read_addr_full_n(mat_B_ch_0_read_addr__full_n),
    .B_read_addr_write(mat_B_ch_0_read_addr__write),
    .B_read_data_s_dout({1'b0, mat_B_ch_0_read_data__dout}),
    .B_read_data_peek_dout({1'b0, mat_B_ch_0_read_data__dout}),
    .B_read_data_s_empty_n(mat_B_ch_0_read_data__empty_n),
    .B_read_data_peek_empty_n(mat_B_ch_0_read_data__empty_n),
    .B_read_data_s_read(mat_B_ch_0_read_data__read),
    .B_read_data_peek_read(),
    .B_write_addr_din(mat_B_ch_0_write_addr__din),
    .B_write_addr_full_n(mat_B_ch_0_write_addr__full_n),
    .B_write_addr_write(mat_B_ch_0_write_addr__write),
    .B_write_data_din(mat_B_ch_0_write_data__din),
    .B_write_data_full_n(mat_B_ch_0_write_data__full_n),
    .B_write_data_write(mat_B_ch_0_write_data__write),
    .B_write_resp_s_dout({1'b0, mat_B_ch_0_write_resp__dout}),
    .B_write_resp_peek_dout({1'b0, mat_B_ch_0_write_resp__dout}),
    .B_write_resp_s_empty_n(mat_B_ch_0_write_resp__empty_n),
    .B_write_resp_peek_empty_n(mat_B_ch_0_write_resp__empty_n),
    .B_write_resp_s_read(mat_B_ch_0_write_resp__read),
    .B_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) read_B
  read_B_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_B_1__ap_start),
    .ap_done(read_B_1__ap_done),
    .ap_idle(read_B_1__ap_idle),
    .ap_ready(read_B_1__ap_ready),
    .K(read_B_1___K__q0),
    .P_N(read_B_1___P_N__q0),
    .fifo_B_din(fifo_B_pe_Sextans_1__din),
    .fifo_B_full_n(fifo_B_pe_Sextans_1__full_n),
    .fifo_B_write(fifo_B_pe_Sextans_1__write),
    .B_read_addr_din(mat_B_ch_1_read_addr__din),
    .B_read_addr_full_n(mat_B_ch_1_read_addr__full_n),
    .B_read_addr_write(mat_B_ch_1_read_addr__write),
    .B_read_data_s_dout({1'b0, mat_B_ch_1_read_data__dout}),
    .B_read_data_peek_dout({1'b0, mat_B_ch_1_read_data__dout}),
    .B_read_data_s_empty_n(mat_B_ch_1_read_data__empty_n),
    .B_read_data_peek_empty_n(mat_B_ch_1_read_data__empty_n),
    .B_read_data_s_read(mat_B_ch_1_read_data__read),
    .B_read_data_peek_read(),
    .B_write_addr_din(mat_B_ch_1_write_addr__din),
    .B_write_addr_full_n(mat_B_ch_1_write_addr__full_n),
    .B_write_addr_write(mat_B_ch_1_write_addr__write),
    .B_write_data_din(mat_B_ch_1_write_data__din),
    .B_write_data_full_n(mat_B_ch_1_write_data__full_n),
    .B_write_data_write(mat_B_ch_1_write_data__write),
    .B_write_resp_s_dout({1'b0, mat_B_ch_1_write_resp__dout}),
    .B_write_resp_peek_dout({1'b0, mat_B_ch_1_write_resp__dout}),
    .B_write_resp_s_empty_n(mat_B_ch_1_write_resp__empty_n),
    .B_write_resp_peek_empty_n(mat_B_ch_1_write_resp__empty_n),
    .B_write_resp_s_read(mat_B_ch_1_write_resp__read),
    .B_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) read_B
  read_B_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_B_2__ap_start),
    .ap_done(read_B_2__ap_done),
    .ap_idle(read_B_2__ap_idle),
    .ap_ready(read_B_2__ap_ready),
    .K(read_B_2___K__q0),
    .P_N(read_B_2___P_N__q0),
    .fifo_B_din(fifo_B_pe_Sextans_2__din),
    .fifo_B_full_n(fifo_B_pe_Sextans_2__full_n),
    .fifo_B_write(fifo_B_pe_Sextans_2__write),
    .B_read_addr_din(mat_B_ch_2_read_addr__din),
    .B_read_addr_full_n(mat_B_ch_2_read_addr__full_n),
    .B_read_addr_write(mat_B_ch_2_read_addr__write),
    .B_read_data_s_dout({1'b0, mat_B_ch_2_read_data__dout}),
    .B_read_data_peek_dout({1'b0, mat_B_ch_2_read_data__dout}),
    .B_read_data_s_empty_n(mat_B_ch_2_read_data__empty_n),
    .B_read_data_peek_empty_n(mat_B_ch_2_read_data__empty_n),
    .B_read_data_s_read(mat_B_ch_2_read_data__read),
    .B_read_data_peek_read(),
    .B_write_addr_din(mat_B_ch_2_write_addr__din),
    .B_write_addr_full_n(mat_B_ch_2_write_addr__full_n),
    .B_write_addr_write(mat_B_ch_2_write_addr__write),
    .B_write_data_din(mat_B_ch_2_write_data__din),
    .B_write_data_full_n(mat_B_ch_2_write_data__full_n),
    .B_write_data_write(mat_B_ch_2_write_data__write),
    .B_write_resp_s_dout({1'b0, mat_B_ch_2_write_resp__dout}),
    .B_write_resp_peek_dout({1'b0, mat_B_ch_2_write_resp__dout}),
    .B_write_resp_s_empty_n(mat_B_ch_2_write_resp__empty_n),
    .B_write_resp_peek_empty_n(mat_B_ch_2_write_resp__empty_n),
    .B_write_resp_s_read(mat_B_ch_2_write_resp__read),
    .B_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) read_B
  read_B_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_B_3__ap_start),
    .ap_done(read_B_3__ap_done),
    .ap_idle(read_B_3__ap_idle),
    .ap_ready(read_B_3__ap_ready),
    .K(read_B_3___K__q0),
    .P_N(read_B_3___P_N__q0),
    .fifo_B_din(fifo_B_pe_Sextans_3__din),
    .fifo_B_full_n(fifo_B_pe_Sextans_3__full_n),
    .fifo_B_write(fifo_B_pe_Sextans_3__write),
    .B_read_addr_din(mat_B_ch_3_read_addr__din),
    .B_read_addr_full_n(mat_B_ch_3_read_addr__full_n),
    .B_read_addr_write(mat_B_ch_3_read_addr__write),
    .B_read_data_s_dout({1'b0, mat_B_ch_3_read_data__dout}),
    .B_read_data_peek_dout({1'b0, mat_B_ch_3_read_data__dout}),
    .B_read_data_s_empty_n(mat_B_ch_3_read_data__empty_n),
    .B_read_data_peek_empty_n(mat_B_ch_3_read_data__empty_n),
    .B_read_data_s_read(mat_B_ch_3_read_data__read),
    .B_read_data_peek_read(),
    .B_write_addr_din(mat_B_ch_3_write_addr__din),
    .B_write_addr_full_n(mat_B_ch_3_write_addr__full_n),
    .B_write_addr_write(mat_B_ch_3_write_addr__write),
    .B_write_data_din(mat_B_ch_3_write_data__din),
    .B_write_data_full_n(mat_B_ch_3_write_data__full_n),
    .B_write_data_write(mat_B_ch_3_write_data__write),
    .B_write_resp_s_dout({1'b0, mat_B_ch_3_write_resp__dout}),
    .B_write_resp_peek_dout({1'b0, mat_B_ch_3_write_resp__dout}),
    .B_write_resp_s_empty_n(mat_B_ch_3_write_resp__empty_n),
    .B_write_resp_peek_empty_n(mat_B_ch_3_write_resp__empty_n),
    .B_write_resp_s_read(mat_B_ch_3_write_resp__read),
    .B_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_0__ap_start),
    .ap_done(read_C_0__ap_done),
    .ap_idle(read_C_0__ap_idle),
    .ap_ready(read_C_0__ap_ready),
    .M(read_C_0___M__q0),
    .P_N(read_C_0___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_0__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_0__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_0__write),
    .C_read_addr_din(mat_C_ch_in_0_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_0_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_0_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_0_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_0_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_0_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_0_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_0_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_0_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_0_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_0_write_addr__write),
    .C_write_data_din(mat_C_ch_in_0_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_0_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_0_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_0_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_0_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_0_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_0_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_0_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_0__din),
    .wrC_inst_full_n(wrC_inst_Sextans_0__full_n),
    .wrC_inst_write(wrC_inst_Sextans_0__write)
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_1__ap_start),
    .ap_done(read_C_1__ap_done),
    .ap_idle(read_C_1__ap_idle),
    .ap_ready(read_C_1__ap_ready),
    .M(read_C_1___M__q0),
    .P_N(read_C_1___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_1__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_1__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_1__write),
    .C_read_addr_din(mat_C_ch_in_1_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_1_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_1_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_1_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_1_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_1_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_1_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_1_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_1_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_1_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_1_write_addr__write),
    .C_write_data_din(mat_C_ch_in_1_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_1_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_1_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_1_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_1_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_1_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_1_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_1_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_1__din),
    .wrC_inst_full_n(wrC_inst_Sextans_1__full_n),
    .wrC_inst_write(wrC_inst_Sextans_1__write)
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_2__ap_start),
    .ap_done(read_C_2__ap_done),
    .ap_idle(read_C_2__ap_idle),
    .ap_ready(read_C_2__ap_ready),
    .M(read_C_2___M__q0),
    .P_N(read_C_2___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_2__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_2__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_2__write),
    .C_read_addr_din(mat_C_ch_in_2_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_2_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_2_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_2_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_2_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_2_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_2_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_2_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_2_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_2_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_2_write_addr__write),
    .C_write_data_din(mat_C_ch_in_2_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_2_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_2_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_2_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_2_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_2_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_2_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_2_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_2__din),
    .wrC_inst_full_n(wrC_inst_Sextans_2__full_n),
    .wrC_inst_write(wrC_inst_Sextans_2__write)
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_3__ap_start),
    .ap_done(read_C_3__ap_done),
    .ap_idle(read_C_3__ap_idle),
    .ap_ready(read_C_3__ap_ready),
    .M(read_C_3___M__q0),
    .P_N(read_C_3___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_3__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_3__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_3__write),
    .C_read_addr_din(mat_C_ch_in_3_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_3_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_3_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_3_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_3_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_3_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_3_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_3_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_3_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_3_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_3_write_addr__write),
    .C_write_data_din(mat_C_ch_in_3_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_3_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_3_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_3_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_3_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_3_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_3_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_3_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_3__din),
    .wrC_inst_full_n(wrC_inst_Sextans_3__full_n),
    .wrC_inst_write(wrC_inst_Sextans_3__write)
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_4__ap_start),
    .ap_done(read_C_4__ap_done),
    .ap_idle(read_C_4__ap_idle),
    .ap_ready(read_C_4__ap_ready),
    .M(read_C_4___M__q0),
    .P_N(read_C_4___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_4__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_4__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_4__write),
    .C_read_addr_din(mat_C_ch_in_4_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_4_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_4_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_4_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_4_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_4_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_4_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_4_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_4_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_4_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_4_write_addr__write),
    .C_write_data_din(mat_C_ch_in_4_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_4_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_4_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_4_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_4_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_4_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_4_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_4_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_4__din),
    .wrC_inst_full_n(wrC_inst_Sextans_4__full_n),
    .wrC_inst_write(wrC_inst_Sextans_4__write)
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_5__ap_start),
    .ap_done(read_C_5__ap_done),
    .ap_idle(read_C_5__ap_idle),
    .ap_ready(read_C_5__ap_ready),
    .M(read_C_5___M__q0),
    .P_N(read_C_5___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_5__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_5__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_5__write),
    .C_read_addr_din(mat_C_ch_in_5_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_5_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_5_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_5_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_5_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_5_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_5_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_5_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_5_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_5_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_5_write_addr__write),
    .C_write_data_din(mat_C_ch_in_5_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_5_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_5_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_5_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_5_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_5_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_5_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_5_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_5__din),
    .wrC_inst_full_n(wrC_inst_Sextans_5__full_n),
    .wrC_inst_write(wrC_inst_Sextans_5__write)
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_6__ap_start),
    .ap_done(read_C_6__ap_done),
    .ap_idle(read_C_6__ap_idle),
    .ap_ready(read_C_6__ap_ready),
    .M(read_C_6___M__q0),
    .P_N(read_C_6___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_6__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_6__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_6__write),
    .C_read_addr_din(mat_C_ch_in_6_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_6_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_6_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_6_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_6_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_6_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_6_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_6_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_6_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_6_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_6_write_addr__write),
    .C_write_data_din(mat_C_ch_in_6_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_6_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_6_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_6_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_6_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_6_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_6_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_6_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_6__din),
    .wrC_inst_full_n(wrC_inst_Sextans_6__full_n),
    .wrC_inst_write(wrC_inst_Sextans_6__write)
  );


  (* keep_hierarchy = "yes" *) read_C
  read_C_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_C_7__ap_start),
    .ap_done(read_C_7__ap_done),
    .ap_idle(read_C_7__ap_idle),
    .ap_ready(read_C_7__ap_ready),
    .M(read_C_7___M__q0),
    .P_N(read_C_7___P_N__q0),
    .fifo_C_din(fifo_C_read_in_Sextans_7__din),
    .fifo_C_full_n(fifo_C_read_in_Sextans_7__full_n),
    .fifo_C_write(fifo_C_read_in_Sextans_7__write),
    .C_read_addr_din(mat_C_ch_in_7_read_addr__din),
    .C_read_addr_full_n(mat_C_ch_in_7_read_addr__full_n),
    .C_read_addr_write(mat_C_ch_in_7_read_addr__write),
    .C_read_data_s_dout({1'b0, mat_C_ch_in_7_read_data__dout}),
    .C_read_data_peek_dout({1'b0, mat_C_ch_in_7_read_data__dout}),
    .C_read_data_s_empty_n(mat_C_ch_in_7_read_data__empty_n),
    .C_read_data_peek_empty_n(mat_C_ch_in_7_read_data__empty_n),
    .C_read_data_s_read(mat_C_ch_in_7_read_data__read),
    .C_read_data_peek_read(),
    .C_write_addr_din(mat_C_ch_in_7_write_addr__din),
    .C_write_addr_full_n(mat_C_ch_in_7_write_addr__full_n),
    .C_write_addr_write(mat_C_ch_in_7_write_addr__write),
    .C_write_data_din(mat_C_ch_in_7_write_data__din),
    .C_write_data_full_n(mat_C_ch_in_7_write_data__full_n),
    .C_write_data_write(mat_C_ch_in_7_write_data__write),
    .C_write_resp_s_dout({1'b0, mat_C_ch_in_7_write_resp__dout}),
    .C_write_resp_peek_dout({1'b0, mat_C_ch_in_7_write_resp__dout}),
    .C_write_resp_s_empty_n(mat_C_ch_in_7_write_resp__empty_n),
    .C_write_resp_peek_empty_n(mat_C_ch_in_7_write_resp__empty_n),
    .C_write_resp_s_read(mat_C_ch_in_7_write_resp__read),
    .C_write_resp_peek_read(),
    .wrC_inst_din(wrC_inst_Sextans_7__din),
    .wrC_inst_full_n(wrC_inst_Sextans_7__full_n),
    .wrC_inst_write(wrC_inst_Sextans_7__write)
  );


  (* keep_hierarchy = "yes" *) read_edge_list_ptr
  read_edge_list_ptr_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(read_edge_list_ptr_0__ap_start),
    .ap_done(read_edge_list_ptr_0__ap_done),
    .ap_idle(read_edge_list_ptr_0__ap_idle),
    .ap_ready(read_edge_list_ptr_0__ap_ready),
    .K(read_edge_list_ptr_0___K__q0),
    .M(read_edge_list_ptr_0___M__q0),
    .num_ite(read_edge_list_ptr_0___NUM_ITE__q0),
    .PE_inst_din(PE_inst_Sextans_0__din),
    .PE_inst_full_n(PE_inst_Sextans_0__full_n),
    .PE_inst_write(PE_inst_Sextans_0__write),
    .P_N(read_edge_list_ptr_0___P_N__q0),
    .edge_list_ptr_read_addr_din(edge_list_ptr_read_addr__din),
    .edge_list_ptr_read_addr_full_n(edge_list_ptr_read_addr__full_n),
    .edge_list_ptr_read_addr_write(edge_list_ptr_read_addr__write),
    .edge_list_ptr_read_data_s_dout({1'b0, edge_list_ptr_read_data__dout}),
    .edge_list_ptr_read_data_peek_dout({1'b0, edge_list_ptr_read_data__dout}),
    .edge_list_ptr_read_data_s_empty_n(edge_list_ptr_read_data__empty_n),
    .edge_list_ptr_read_data_peek_empty_n(edge_list_ptr_read_data__empty_n),
    .edge_list_ptr_read_data_s_read(edge_list_ptr_read_data__read),
    .edge_list_ptr_read_data_peek_read(),
    .edge_list_ptr_write_addr_din(edge_list_ptr_write_addr__din),
    .edge_list_ptr_write_addr_full_n(edge_list_ptr_write_addr__full_n),
    .edge_list_ptr_write_addr_write(edge_list_ptr_write_addr__write),
    .edge_list_ptr_write_data_din(edge_list_ptr_write_data__din),
    .edge_list_ptr_write_data_full_n(edge_list_ptr_write_data__full_n),
    .edge_list_ptr_write_data_write(edge_list_ptr_write_data__write),
    .edge_list_ptr_write_resp_s_dout({1'b0, edge_list_ptr_write_resp__dout}),
    .edge_list_ptr_write_resp_peek_dout({1'b0, edge_list_ptr_write_resp__dout}),
    .edge_list_ptr_write_resp_s_empty_n(edge_list_ptr_write_resp__empty_n),
    .edge_list_ptr_write_resp_peek_empty_n(edge_list_ptr_write_resp__empty_n),
    .edge_list_ptr_write_resp_s_read(edge_list_ptr_write_resp__read),
    .edge_list_ptr_write_resp_peek_read(),
    .fifo_edge_list_ptr_din(fifo_edge_list_ptr_Sextans_0__din),
    .fifo_edge_list_ptr_full_n(fifo_edge_list_ptr_Sextans_0__full_n),
    .fifo_edge_list_ptr_write(fifo_edge_list_ptr_Sextans_0__write)
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_0__ap_start),
    .ap_done(write_C_0__ap_done),
    .ap_idle(write_C_0__ap_idle),
    .ap_ready(write_C_0__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_0__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_0__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_0__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_0__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_0__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_0_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_0_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_0_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_0_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_0_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_0_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_0_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_0_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_0_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_0_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_0_write_addr__write),
    .C_out_write_data_din(mat_C_ch_0_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_0_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_0_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_0_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_0_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_0_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_0_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_0_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_0__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_0__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_0__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_0__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_0__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_1__ap_start),
    .ap_done(write_C_1__ap_done),
    .ap_idle(write_C_1__ap_idle),
    .ap_ready(write_C_1__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_1__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_1__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_1__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_1__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_1__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_1_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_1_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_1_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_1_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_1_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_1_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_1_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_1_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_1_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_1_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_1_write_addr__write),
    .C_out_write_data_din(mat_C_ch_1_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_1_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_1_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_1_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_1_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_1_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_1_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_1_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_1__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_1__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_1__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_1__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_1__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_2__ap_start),
    .ap_done(write_C_2__ap_done),
    .ap_idle(write_C_2__ap_idle),
    .ap_ready(write_C_2__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_2__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_2__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_2__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_2__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_2__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_2_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_2_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_2_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_2_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_2_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_2_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_2_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_2_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_2_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_2_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_2_write_addr__write),
    .C_out_write_data_din(mat_C_ch_2_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_2_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_2_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_2_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_2_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_2_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_2_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_2_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_2__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_2__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_2__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_2__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_2__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_3__ap_start),
    .ap_done(write_C_3__ap_done),
    .ap_idle(write_C_3__ap_idle),
    .ap_ready(write_C_3__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_3__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_3__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_3__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_3__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_3__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_3_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_3_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_3_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_3_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_3_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_3_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_3_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_3_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_3_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_3_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_3_write_addr__write),
    .C_out_write_data_din(mat_C_ch_3_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_3_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_3_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_3_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_3_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_3_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_3_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_3_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_3__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_3__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_3__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_3__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_3__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_4__ap_start),
    .ap_done(write_C_4__ap_done),
    .ap_idle(write_C_4__ap_idle),
    .ap_ready(write_C_4__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_4__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_4__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_4__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_4__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_4__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_4_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_4_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_4_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_4_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_4_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_4_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_4_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_4_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_4_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_4_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_4_write_addr__write),
    .C_out_write_data_din(mat_C_ch_4_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_4_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_4_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_4_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_4_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_4_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_4_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_4_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_4__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_4__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_4__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_4__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_4__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_5__ap_start),
    .ap_done(write_C_5__ap_done),
    .ap_idle(write_C_5__ap_idle),
    .ap_ready(write_C_5__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_5__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_5__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_5__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_5__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_5__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_5_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_5_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_5_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_5_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_5_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_5_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_5_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_5_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_5_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_5_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_5_write_addr__write),
    .C_out_write_data_din(mat_C_ch_5_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_5_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_5_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_5_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_5_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_5_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_5_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_5_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_5__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_5__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_5__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_5__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_5__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_6__ap_start),
    .ap_done(write_C_6__ap_done),
    .ap_idle(write_C_6__ap_idle),
    .ap_ready(write_C_6__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_6__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_6__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_6__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_6__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_6__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_6_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_6_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_6_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_6_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_6_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_6_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_6_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_6_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_6_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_6_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_6_write_addr__write),
    .C_out_write_data_din(mat_C_ch_6_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_6_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_6_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_6_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_6_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_6_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_6_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_6_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_6__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_6__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_6__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_6__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_6__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) write_C
  write_C_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(write_C_7__ap_start),
    .ap_done(write_C_7__ap_done),
    .ap_idle(write_C_7__ap_idle),
    .ap_ready(write_C_7__ap_ready),
    .fifo_C_s_dout(fifo_C_ch_Sextans_7__dout),
    .fifo_C_peek_dout(fifo_C_ch_Sextans_7__dout),
    .fifo_C_s_empty_n(fifo_C_ch_Sextans_7__empty_n),
    .fifo_C_peek_empty_n(fifo_C_ch_Sextans_7__empty_n),
    .fifo_C_s_read(fifo_C_ch_Sextans_7__read),
    .fifo_C_peek_read(),
    .C_out_read_addr_din(mat_C_ch_7_read_addr__din),
    .C_out_read_addr_full_n(mat_C_ch_7_read_addr__full_n),
    .C_out_read_addr_write(mat_C_ch_7_read_addr__write),
    .C_out_read_data_s_dout({1'b0, mat_C_ch_7_read_data__dout}),
    .C_out_read_data_peek_dout({1'b0, mat_C_ch_7_read_data__dout}),
    .C_out_read_data_s_empty_n(mat_C_ch_7_read_data__empty_n),
    .C_out_read_data_peek_empty_n(mat_C_ch_7_read_data__empty_n),
    .C_out_read_data_s_read(mat_C_ch_7_read_data__read),
    .C_out_read_data_peek_read(),
    .C_out_write_addr_din(mat_C_ch_7_write_addr__din),
    .C_out_write_addr_full_n(mat_C_ch_7_write_addr__full_n),
    .C_out_write_addr_write(mat_C_ch_7_write_addr__write),
    .C_out_write_data_din(mat_C_ch_7_write_data__din),
    .C_out_write_data_full_n(mat_C_ch_7_write_data__full_n),
    .C_out_write_data_write(mat_C_ch_7_write_data__write),
    .C_out_write_resp_s_dout({1'b0, mat_C_ch_7_write_resp__dout}),
    .C_out_write_resp_peek_dout({1'b0, mat_C_ch_7_write_resp__dout}),
    .C_out_write_resp_s_empty_n(mat_C_ch_7_write_resp__empty_n),
    .C_out_write_resp_peek_empty_n(mat_C_ch_7_write_resp__empty_n),
    .C_out_write_resp_s_read(mat_C_ch_7_write_resp__read),
    .C_out_write_resp_peek_read(),
    .wrC_inst_s_dout(wrC_inst_Sextans_7__dout),
    .wrC_inst_peek_dout(wrC_inst_Sextans_7__dout),
    .wrC_inst_s_empty_n(wrC_inst_Sextans_7__empty_n),
    .wrC_inst_peek_empty_n(wrC_inst_Sextans_7__empty_n),
    .wrC_inst_s_read(wrC_inst_Sextans_7__read),
    .wrC_inst_peek_read()
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_0___edge_list_ch_0__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_0_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_0_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_0_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_0_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_0_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_0_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_0_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_0_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_0_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_0_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_0_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_0_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_0_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_0_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_0_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_0_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_0_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_0_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_0_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_0_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_0_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_0_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_0_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_0_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_0_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_0_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_0_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_0_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_0_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_0_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_0_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_0_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_0_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_0_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_0_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_0_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_0_WVALID),
    .read_addr_din(edge_list_ch_0_read_addr__din),
    .read_addr_full_n(edge_list_ch_0_read_addr__full_n),
    .read_addr_write(edge_list_ch_0_read_addr__write),
    .read_data_dout(edge_list_ch_0_read_data__dout),
    .read_data_empty_n(edge_list_ch_0_read_data__empty_n),
    .read_data_read(edge_list_ch_0_read_data__read),
    .write_addr_din(edge_list_ch_0_write_addr__din),
    .write_addr_full_n(edge_list_ch_0_write_addr__full_n),
    .write_addr_write(edge_list_ch_0_write_addr__write),
    .write_data_din(edge_list_ch_0_write_data__din),
    .write_data_full_n(edge_list_ch_0_write_data__full_n),
    .write_data_write(edge_list_ch_0_write_data__write),
    .write_resp_dout(edge_list_ch_0_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_0_write_resp__empty_n),
    .write_resp_read(edge_list_ch_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_1___edge_list_ch_1__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_1_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_1_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_1_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_1_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_1_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_1_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_1_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_1_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_1_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_1_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_1_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_1_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_1_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_1_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_1_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_1_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_1_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_1_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_1_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_1_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_1_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_1_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_1_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_1_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_1_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_1_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_1_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_1_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_1_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_1_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_1_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_1_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_1_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_1_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_1_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_1_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_1_WVALID),
    .read_addr_din(edge_list_ch_1_read_addr__din),
    .read_addr_full_n(edge_list_ch_1_read_addr__full_n),
    .read_addr_write(edge_list_ch_1_read_addr__write),
    .read_data_dout(edge_list_ch_1_read_data__dout),
    .read_data_empty_n(edge_list_ch_1_read_data__empty_n),
    .read_data_read(edge_list_ch_1_read_data__read),
    .write_addr_din(edge_list_ch_1_write_addr__din),
    .write_addr_full_n(edge_list_ch_1_write_addr__full_n),
    .write_addr_write(edge_list_ch_1_write_addr__write),
    .write_data_din(edge_list_ch_1_write_data__din),
    .write_data_full_n(edge_list_ch_1_write_data__full_n),
    .write_data_write(edge_list_ch_1_write_data__write),
    .write_resp_dout(edge_list_ch_1_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_1_write_resp__empty_n),
    .write_resp_read(edge_list_ch_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_2___edge_list_ch_2__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_2_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_2_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_2_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_2_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_2_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_2_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_2_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_2_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_2_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_2_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_2_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_2_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_2_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_2_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_2_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_2_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_2_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_2_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_2_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_2_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_2_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_2_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_2_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_2_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_2_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_2_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_2_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_2_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_2_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_2_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_2_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_2_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_2_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_2_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_2_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_2_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_2_WVALID),
    .read_addr_din(edge_list_ch_2_read_addr__din),
    .read_addr_full_n(edge_list_ch_2_read_addr__full_n),
    .read_addr_write(edge_list_ch_2_read_addr__write),
    .read_data_dout(edge_list_ch_2_read_data__dout),
    .read_data_empty_n(edge_list_ch_2_read_data__empty_n),
    .read_data_read(edge_list_ch_2_read_data__read),
    .write_addr_din(edge_list_ch_2_write_addr__din),
    .write_addr_full_n(edge_list_ch_2_write_addr__full_n),
    .write_addr_write(edge_list_ch_2_write_addr__write),
    .write_data_din(edge_list_ch_2_write_data__din),
    .write_data_full_n(edge_list_ch_2_write_data__full_n),
    .write_data_write(edge_list_ch_2_write_data__write),
    .write_resp_dout(edge_list_ch_2_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_2_write_resp__empty_n),
    .write_resp_read(edge_list_ch_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_3___edge_list_ch_3__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_3_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_3_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_3_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_3_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_3_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_3_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_3_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_3_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_3_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_3_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_3_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_3_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_3_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_3_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_3_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_3_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_3_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_3_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_3_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_3_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_3_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_3_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_3_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_3_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_3_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_3_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_3_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_3_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_3_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_3_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_3_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_3_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_3_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_3_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_3_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_3_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_3_WVALID),
    .read_addr_din(edge_list_ch_3_read_addr__din),
    .read_addr_full_n(edge_list_ch_3_read_addr__full_n),
    .read_addr_write(edge_list_ch_3_read_addr__write),
    .read_data_dout(edge_list_ch_3_read_data__dout),
    .read_data_empty_n(edge_list_ch_3_read_data__empty_n),
    .read_data_read(edge_list_ch_3_read_data__read),
    .write_addr_din(edge_list_ch_3_write_addr__din),
    .write_addr_full_n(edge_list_ch_3_write_addr__full_n),
    .write_addr_write(edge_list_ch_3_write_addr__write),
    .write_data_din(edge_list_ch_3_write_data__din),
    .write_data_full_n(edge_list_ch_3_write_data__full_n),
    .write_data_write(edge_list_ch_3_write_data__write),
    .write_resp_dout(edge_list_ch_3_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_3_write_resp__empty_n),
    .write_resp_read(edge_list_ch_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_4__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_4___edge_list_ch_4__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_4_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_4_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_4_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_4_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_4_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_4_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_4_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_4_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_4_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_4_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_4_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_4_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_4_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_4_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_4_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_4_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_4_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_4_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_4_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_4_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_4_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_4_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_4_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_4_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_4_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_4_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_4_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_4_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_4_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_4_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_4_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_4_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_4_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_4_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_4_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_4_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_4_WVALID),
    .read_addr_din(edge_list_ch_4_read_addr__din),
    .read_addr_full_n(edge_list_ch_4_read_addr__full_n),
    .read_addr_write(edge_list_ch_4_read_addr__write),
    .read_data_dout(edge_list_ch_4_read_data__dout),
    .read_data_empty_n(edge_list_ch_4_read_data__empty_n),
    .read_data_read(edge_list_ch_4_read_data__read),
    .write_addr_din(edge_list_ch_4_write_addr__din),
    .write_addr_full_n(edge_list_ch_4_write_addr__full_n),
    .write_addr_write(edge_list_ch_4_write_addr__write),
    .write_data_din(edge_list_ch_4_write_data__din),
    .write_data_full_n(edge_list_ch_4_write_data__full_n),
    .write_data_write(edge_list_ch_4_write_data__write),
    .write_resp_dout(edge_list_ch_4_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_4_write_resp__empty_n),
    .write_resp_read(edge_list_ch_4_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_5__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_5___edge_list_ch_5__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_5_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_5_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_5_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_5_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_5_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_5_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_5_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_5_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_5_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_5_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_5_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_5_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_5_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_5_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_5_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_5_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_5_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_5_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_5_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_5_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_5_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_5_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_5_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_5_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_5_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_5_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_5_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_5_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_5_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_5_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_5_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_5_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_5_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_5_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_5_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_5_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_5_WVALID),
    .read_addr_din(edge_list_ch_5_read_addr__din),
    .read_addr_full_n(edge_list_ch_5_read_addr__full_n),
    .read_addr_write(edge_list_ch_5_read_addr__write),
    .read_data_dout(edge_list_ch_5_read_data__dout),
    .read_data_empty_n(edge_list_ch_5_read_data__empty_n),
    .read_data_read(edge_list_ch_5_read_data__read),
    .write_addr_din(edge_list_ch_5_write_addr__din),
    .write_addr_full_n(edge_list_ch_5_write_addr__full_n),
    .write_addr_write(edge_list_ch_5_write_addr__write),
    .write_data_din(edge_list_ch_5_write_data__din),
    .write_data_full_n(edge_list_ch_5_write_data__full_n),
    .write_data_write(edge_list_ch_5_write_data__write),
    .write_resp_dout(edge_list_ch_5_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_5_write_resp__empty_n),
    .write_resp_read(edge_list_ch_5_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_6__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_6___edge_list_ch_6__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_6_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_6_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_6_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_6_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_6_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_6_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_6_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_6_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_6_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_6_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_6_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_6_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_6_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_6_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_6_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_6_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_6_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_6_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_6_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_6_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_6_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_6_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_6_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_6_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_6_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_6_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_6_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_6_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_6_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_6_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_6_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_6_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_6_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_6_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_6_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_6_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_6_WVALID),
    .read_addr_din(edge_list_ch_6_read_addr__din),
    .read_addr_full_n(edge_list_ch_6_read_addr__full_n),
    .read_addr_write(edge_list_ch_6_read_addr__write),
    .read_data_dout(edge_list_ch_6_read_data__dout),
    .read_data_empty_n(edge_list_ch_6_read_data__empty_n),
    .read_data_read(edge_list_ch_6_read_data__read),
    .write_addr_din(edge_list_ch_6_write_addr__din),
    .write_addr_full_n(edge_list_ch_6_write_addr__full_n),
    .write_addr_write(edge_list_ch_6_write_addr__write),
    .write_data_din(edge_list_ch_6_write_data__din),
    .write_data_full_n(edge_list_ch_6_write_data__full_n),
    .write_data_write(edge_list_ch_6_write_data__write),
    .write_resp_dout(edge_list_ch_6_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_6_write_resp__empty_n),
    .write_resp_read(edge_list_ch_6_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  edge_list_ch_7__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_A_7___edge_list_ch_7__q0),
    .m_axi_ARADDR(m_axi_edge_list_ch_7_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ch_7_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ch_7_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ch_7_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ch_7_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ch_7_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ch_7_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ch_7_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ch_7_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ch_7_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ch_7_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ch_7_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ch_7_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ch_7_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ch_7_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ch_7_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ch_7_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ch_7_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ch_7_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ch_7_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ch_7_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ch_7_AWVALID),
    .m_axi_BID(m_axi_edge_list_ch_7_BID),
    .m_axi_BREADY(m_axi_edge_list_ch_7_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ch_7_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ch_7_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ch_7_RDATA),
    .m_axi_RID(m_axi_edge_list_ch_7_RID),
    .m_axi_RLAST(m_axi_edge_list_ch_7_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ch_7_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ch_7_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ch_7_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ch_7_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ch_7_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ch_7_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ch_7_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ch_7_WVALID),
    .read_addr_din(edge_list_ch_7_read_addr__din),
    .read_addr_full_n(edge_list_ch_7_read_addr__full_n),
    .read_addr_write(edge_list_ch_7_read_addr__write),
    .read_data_dout(edge_list_ch_7_read_data__dout),
    .read_data_empty_n(edge_list_ch_7_read_data__empty_n),
    .read_data_read(edge_list_ch_7_read_data__read),
    .write_addr_din(edge_list_ch_7_write_addr__din),
    .write_addr_full_n(edge_list_ch_7_write_addr__full_n),
    .write_addr_write(edge_list_ch_7_write_addr__write),
    .write_data_din(edge_list_ch_7_write_data__din),
    .write_data_full_n(edge_list_ch_7_write_data__full_n),
    .write_data_write(edge_list_ch_7_write_data__write),
    .write_resp_dout(edge_list_ch_7_write_resp__dout),
    .write_resp_empty_n(edge_list_ch_7_write_resp__empty_n),
    .write_resp_read(edge_list_ch_7_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_B_ch_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_B_0___mat_B_ch_0__q0),
    .m_axi_ARADDR(m_axi_mat_B_ch_0_ARADDR),
    .m_axi_ARBURST(m_axi_mat_B_ch_0_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_B_ch_0_ARCACHE),
    .m_axi_ARID(m_axi_mat_B_ch_0_ARID),
    .m_axi_ARLEN(m_axi_mat_B_ch_0_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_B_ch_0_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_B_ch_0_ARPROT),
    .m_axi_ARQOS(m_axi_mat_B_ch_0_ARQOS),
    .m_axi_ARREADY(m_axi_mat_B_ch_0_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_B_ch_0_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_B_ch_0_ARVALID),
    .m_axi_AWADDR(m_axi_mat_B_ch_0_AWADDR),
    .m_axi_AWBURST(m_axi_mat_B_ch_0_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_B_ch_0_AWCACHE),
    .m_axi_AWID(m_axi_mat_B_ch_0_AWID),
    .m_axi_AWLEN(m_axi_mat_B_ch_0_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_B_ch_0_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_B_ch_0_AWPROT),
    .m_axi_AWQOS(m_axi_mat_B_ch_0_AWQOS),
    .m_axi_AWREADY(m_axi_mat_B_ch_0_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_B_ch_0_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_B_ch_0_AWVALID),
    .m_axi_BID(m_axi_mat_B_ch_0_BID),
    .m_axi_BREADY(m_axi_mat_B_ch_0_BREADY),
    .m_axi_BRESP(m_axi_mat_B_ch_0_BRESP),
    .m_axi_BVALID(m_axi_mat_B_ch_0_BVALID),
    .m_axi_RDATA(m_axi_mat_B_ch_0_RDATA),
    .m_axi_RID(m_axi_mat_B_ch_0_RID),
    .m_axi_RLAST(m_axi_mat_B_ch_0_RLAST),
    .m_axi_RREADY(m_axi_mat_B_ch_0_RREADY),
    .m_axi_RRESP(m_axi_mat_B_ch_0_RRESP),
    .m_axi_RVALID(m_axi_mat_B_ch_0_RVALID),
    .m_axi_WDATA(m_axi_mat_B_ch_0_WDATA),
    .m_axi_WLAST(m_axi_mat_B_ch_0_WLAST),
    .m_axi_WREADY(m_axi_mat_B_ch_0_WREADY),
    .m_axi_WSTRB(m_axi_mat_B_ch_0_WSTRB),
    .m_axi_WVALID(m_axi_mat_B_ch_0_WVALID),
    .read_addr_din(mat_B_ch_0_read_addr__din),
    .read_addr_full_n(mat_B_ch_0_read_addr__full_n),
    .read_addr_write(mat_B_ch_0_read_addr__write),
    .read_data_dout(mat_B_ch_0_read_data__dout),
    .read_data_empty_n(mat_B_ch_0_read_data__empty_n),
    .read_data_read(mat_B_ch_0_read_data__read),
    .write_addr_din(mat_B_ch_0_write_addr__din),
    .write_addr_full_n(mat_B_ch_0_write_addr__full_n),
    .write_addr_write(mat_B_ch_0_write_addr__write),
    .write_data_din(mat_B_ch_0_write_data__din),
    .write_data_full_n(mat_B_ch_0_write_data__full_n),
    .write_data_write(mat_B_ch_0_write_data__write),
    .write_resp_dout(mat_B_ch_0_write_resp__dout),
    .write_resp_empty_n(mat_B_ch_0_write_resp__empty_n),
    .write_resp_read(mat_B_ch_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_B_ch_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_B_1___mat_B_ch_1__q0),
    .m_axi_ARADDR(m_axi_mat_B_ch_1_ARADDR),
    .m_axi_ARBURST(m_axi_mat_B_ch_1_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_B_ch_1_ARCACHE),
    .m_axi_ARID(m_axi_mat_B_ch_1_ARID),
    .m_axi_ARLEN(m_axi_mat_B_ch_1_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_B_ch_1_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_B_ch_1_ARPROT),
    .m_axi_ARQOS(m_axi_mat_B_ch_1_ARQOS),
    .m_axi_ARREADY(m_axi_mat_B_ch_1_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_B_ch_1_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_B_ch_1_ARVALID),
    .m_axi_AWADDR(m_axi_mat_B_ch_1_AWADDR),
    .m_axi_AWBURST(m_axi_mat_B_ch_1_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_B_ch_1_AWCACHE),
    .m_axi_AWID(m_axi_mat_B_ch_1_AWID),
    .m_axi_AWLEN(m_axi_mat_B_ch_1_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_B_ch_1_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_B_ch_1_AWPROT),
    .m_axi_AWQOS(m_axi_mat_B_ch_1_AWQOS),
    .m_axi_AWREADY(m_axi_mat_B_ch_1_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_B_ch_1_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_B_ch_1_AWVALID),
    .m_axi_BID(m_axi_mat_B_ch_1_BID),
    .m_axi_BREADY(m_axi_mat_B_ch_1_BREADY),
    .m_axi_BRESP(m_axi_mat_B_ch_1_BRESP),
    .m_axi_BVALID(m_axi_mat_B_ch_1_BVALID),
    .m_axi_RDATA(m_axi_mat_B_ch_1_RDATA),
    .m_axi_RID(m_axi_mat_B_ch_1_RID),
    .m_axi_RLAST(m_axi_mat_B_ch_1_RLAST),
    .m_axi_RREADY(m_axi_mat_B_ch_1_RREADY),
    .m_axi_RRESP(m_axi_mat_B_ch_1_RRESP),
    .m_axi_RVALID(m_axi_mat_B_ch_1_RVALID),
    .m_axi_WDATA(m_axi_mat_B_ch_1_WDATA),
    .m_axi_WLAST(m_axi_mat_B_ch_1_WLAST),
    .m_axi_WREADY(m_axi_mat_B_ch_1_WREADY),
    .m_axi_WSTRB(m_axi_mat_B_ch_1_WSTRB),
    .m_axi_WVALID(m_axi_mat_B_ch_1_WVALID),
    .read_addr_din(mat_B_ch_1_read_addr__din),
    .read_addr_full_n(mat_B_ch_1_read_addr__full_n),
    .read_addr_write(mat_B_ch_1_read_addr__write),
    .read_data_dout(mat_B_ch_1_read_data__dout),
    .read_data_empty_n(mat_B_ch_1_read_data__empty_n),
    .read_data_read(mat_B_ch_1_read_data__read),
    .write_addr_din(mat_B_ch_1_write_addr__din),
    .write_addr_full_n(mat_B_ch_1_write_addr__full_n),
    .write_addr_write(mat_B_ch_1_write_addr__write),
    .write_data_din(mat_B_ch_1_write_data__din),
    .write_data_full_n(mat_B_ch_1_write_data__full_n),
    .write_data_write(mat_B_ch_1_write_data__write),
    .write_resp_dout(mat_B_ch_1_write_resp__dout),
    .write_resp_empty_n(mat_B_ch_1_write_resp__empty_n),
    .write_resp_read(mat_B_ch_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_B_ch_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_B_2___mat_B_ch_2__q0),
    .m_axi_ARADDR(m_axi_mat_B_ch_2_ARADDR),
    .m_axi_ARBURST(m_axi_mat_B_ch_2_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_B_ch_2_ARCACHE),
    .m_axi_ARID(m_axi_mat_B_ch_2_ARID),
    .m_axi_ARLEN(m_axi_mat_B_ch_2_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_B_ch_2_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_B_ch_2_ARPROT),
    .m_axi_ARQOS(m_axi_mat_B_ch_2_ARQOS),
    .m_axi_ARREADY(m_axi_mat_B_ch_2_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_B_ch_2_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_B_ch_2_ARVALID),
    .m_axi_AWADDR(m_axi_mat_B_ch_2_AWADDR),
    .m_axi_AWBURST(m_axi_mat_B_ch_2_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_B_ch_2_AWCACHE),
    .m_axi_AWID(m_axi_mat_B_ch_2_AWID),
    .m_axi_AWLEN(m_axi_mat_B_ch_2_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_B_ch_2_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_B_ch_2_AWPROT),
    .m_axi_AWQOS(m_axi_mat_B_ch_2_AWQOS),
    .m_axi_AWREADY(m_axi_mat_B_ch_2_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_B_ch_2_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_B_ch_2_AWVALID),
    .m_axi_BID(m_axi_mat_B_ch_2_BID),
    .m_axi_BREADY(m_axi_mat_B_ch_2_BREADY),
    .m_axi_BRESP(m_axi_mat_B_ch_2_BRESP),
    .m_axi_BVALID(m_axi_mat_B_ch_2_BVALID),
    .m_axi_RDATA(m_axi_mat_B_ch_2_RDATA),
    .m_axi_RID(m_axi_mat_B_ch_2_RID),
    .m_axi_RLAST(m_axi_mat_B_ch_2_RLAST),
    .m_axi_RREADY(m_axi_mat_B_ch_2_RREADY),
    .m_axi_RRESP(m_axi_mat_B_ch_2_RRESP),
    .m_axi_RVALID(m_axi_mat_B_ch_2_RVALID),
    .m_axi_WDATA(m_axi_mat_B_ch_2_WDATA),
    .m_axi_WLAST(m_axi_mat_B_ch_2_WLAST),
    .m_axi_WREADY(m_axi_mat_B_ch_2_WREADY),
    .m_axi_WSTRB(m_axi_mat_B_ch_2_WSTRB),
    .m_axi_WVALID(m_axi_mat_B_ch_2_WVALID),
    .read_addr_din(mat_B_ch_2_read_addr__din),
    .read_addr_full_n(mat_B_ch_2_read_addr__full_n),
    .read_addr_write(mat_B_ch_2_read_addr__write),
    .read_data_dout(mat_B_ch_2_read_data__dout),
    .read_data_empty_n(mat_B_ch_2_read_data__empty_n),
    .read_data_read(mat_B_ch_2_read_data__read),
    .write_addr_din(mat_B_ch_2_write_addr__din),
    .write_addr_full_n(mat_B_ch_2_write_addr__full_n),
    .write_addr_write(mat_B_ch_2_write_addr__write),
    .write_data_din(mat_B_ch_2_write_data__din),
    .write_data_full_n(mat_B_ch_2_write_data__full_n),
    .write_data_write(mat_B_ch_2_write_data__write),
    .write_resp_dout(mat_B_ch_2_write_resp__dout),
    .write_resp_empty_n(mat_B_ch_2_write_resp__empty_n),
    .write_resp_read(mat_B_ch_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_B_ch_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_B_3___mat_B_ch_3__q0),
    .m_axi_ARADDR(m_axi_mat_B_ch_3_ARADDR),
    .m_axi_ARBURST(m_axi_mat_B_ch_3_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_B_ch_3_ARCACHE),
    .m_axi_ARID(m_axi_mat_B_ch_3_ARID),
    .m_axi_ARLEN(m_axi_mat_B_ch_3_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_B_ch_3_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_B_ch_3_ARPROT),
    .m_axi_ARQOS(m_axi_mat_B_ch_3_ARQOS),
    .m_axi_ARREADY(m_axi_mat_B_ch_3_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_B_ch_3_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_B_ch_3_ARVALID),
    .m_axi_AWADDR(m_axi_mat_B_ch_3_AWADDR),
    .m_axi_AWBURST(m_axi_mat_B_ch_3_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_B_ch_3_AWCACHE),
    .m_axi_AWID(m_axi_mat_B_ch_3_AWID),
    .m_axi_AWLEN(m_axi_mat_B_ch_3_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_B_ch_3_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_B_ch_3_AWPROT),
    .m_axi_AWQOS(m_axi_mat_B_ch_3_AWQOS),
    .m_axi_AWREADY(m_axi_mat_B_ch_3_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_B_ch_3_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_B_ch_3_AWVALID),
    .m_axi_BID(m_axi_mat_B_ch_3_BID),
    .m_axi_BREADY(m_axi_mat_B_ch_3_BREADY),
    .m_axi_BRESP(m_axi_mat_B_ch_3_BRESP),
    .m_axi_BVALID(m_axi_mat_B_ch_3_BVALID),
    .m_axi_RDATA(m_axi_mat_B_ch_3_RDATA),
    .m_axi_RID(m_axi_mat_B_ch_3_RID),
    .m_axi_RLAST(m_axi_mat_B_ch_3_RLAST),
    .m_axi_RREADY(m_axi_mat_B_ch_3_RREADY),
    .m_axi_RRESP(m_axi_mat_B_ch_3_RRESP),
    .m_axi_RVALID(m_axi_mat_B_ch_3_RVALID),
    .m_axi_WDATA(m_axi_mat_B_ch_3_WDATA),
    .m_axi_WLAST(m_axi_mat_B_ch_3_WLAST),
    .m_axi_WREADY(m_axi_mat_B_ch_3_WREADY),
    .m_axi_WSTRB(m_axi_mat_B_ch_3_WSTRB),
    .m_axi_WVALID(m_axi_mat_B_ch_3_WVALID),
    .read_addr_din(mat_B_ch_3_read_addr__din),
    .read_addr_full_n(mat_B_ch_3_read_addr__full_n),
    .read_addr_write(mat_B_ch_3_read_addr__write),
    .read_data_dout(mat_B_ch_3_read_data__dout),
    .read_data_empty_n(mat_B_ch_3_read_data__empty_n),
    .read_data_read(mat_B_ch_3_read_data__read),
    .write_addr_din(mat_B_ch_3_write_addr__din),
    .write_addr_full_n(mat_B_ch_3_write_addr__full_n),
    .write_addr_write(mat_B_ch_3_write_addr__write),
    .write_data_din(mat_B_ch_3_write_data__din),
    .write_data_full_n(mat_B_ch_3_write_data__full_n),
    .write_data_write(mat_B_ch_3_write_data__write),
    .write_resp_dout(mat_B_ch_3_write_resp__dout),
    .write_resp_empty_n(mat_B_ch_3_write_resp__empty_n),
    .write_resp_read(mat_B_ch_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_0___mat_C_ch_in_0__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_0_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_0_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_0_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_0_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_0_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_0_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_0_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_0_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_0_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_0_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_0_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_0_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_0_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_0_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_0_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_0_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_0_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_0_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_0_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_0_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_0_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_0_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_0_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_0_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_0_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_0_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_0_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_0_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_0_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_0_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_0_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_0_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_0_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_0_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_0_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_0_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_0_WVALID),
    .read_addr_din(mat_C_ch_in_0_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_0_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_0_read_addr__write),
    .read_data_dout(mat_C_ch_in_0_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_0_read_data__empty_n),
    .read_data_read(mat_C_ch_in_0_read_data__read),
    .write_addr_din(mat_C_ch_in_0_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_0_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_0_write_addr__write),
    .write_data_din(mat_C_ch_in_0_write_data__din),
    .write_data_full_n(mat_C_ch_in_0_write_data__full_n),
    .write_data_write(mat_C_ch_in_0_write_data__write),
    .write_resp_dout(mat_C_ch_in_0_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_0_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_1___mat_C_ch_in_1__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_1_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_1_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_1_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_1_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_1_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_1_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_1_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_1_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_1_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_1_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_1_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_1_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_1_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_1_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_1_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_1_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_1_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_1_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_1_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_1_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_1_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_1_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_1_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_1_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_1_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_1_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_1_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_1_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_1_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_1_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_1_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_1_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_1_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_1_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_1_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_1_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_1_WVALID),
    .read_addr_din(mat_C_ch_in_1_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_1_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_1_read_addr__write),
    .read_data_dout(mat_C_ch_in_1_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_1_read_data__empty_n),
    .read_data_read(mat_C_ch_in_1_read_data__read),
    .write_addr_din(mat_C_ch_in_1_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_1_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_1_write_addr__write),
    .write_data_din(mat_C_ch_in_1_write_data__din),
    .write_data_full_n(mat_C_ch_in_1_write_data__full_n),
    .write_data_write(mat_C_ch_in_1_write_data__write),
    .write_resp_dout(mat_C_ch_in_1_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_1_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_2___mat_C_ch_in_2__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_2_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_2_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_2_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_2_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_2_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_2_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_2_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_2_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_2_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_2_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_2_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_2_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_2_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_2_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_2_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_2_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_2_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_2_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_2_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_2_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_2_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_2_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_2_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_2_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_2_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_2_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_2_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_2_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_2_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_2_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_2_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_2_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_2_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_2_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_2_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_2_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_2_WVALID),
    .read_addr_din(mat_C_ch_in_2_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_2_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_2_read_addr__write),
    .read_data_dout(mat_C_ch_in_2_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_2_read_data__empty_n),
    .read_data_read(mat_C_ch_in_2_read_data__read),
    .write_addr_din(mat_C_ch_in_2_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_2_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_2_write_addr__write),
    .write_data_din(mat_C_ch_in_2_write_data__din),
    .write_data_full_n(mat_C_ch_in_2_write_data__full_n),
    .write_data_write(mat_C_ch_in_2_write_data__write),
    .write_resp_dout(mat_C_ch_in_2_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_2_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_3___mat_C_ch_in_3__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_3_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_3_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_3_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_3_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_3_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_3_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_3_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_3_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_3_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_3_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_3_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_3_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_3_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_3_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_3_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_3_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_3_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_3_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_3_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_3_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_3_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_3_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_3_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_3_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_3_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_3_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_3_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_3_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_3_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_3_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_3_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_3_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_3_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_3_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_3_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_3_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_3_WVALID),
    .read_addr_din(mat_C_ch_in_3_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_3_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_3_read_addr__write),
    .read_data_dout(mat_C_ch_in_3_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_3_read_data__empty_n),
    .read_data_read(mat_C_ch_in_3_read_data__read),
    .write_addr_din(mat_C_ch_in_3_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_3_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_3_write_addr__write),
    .write_data_din(mat_C_ch_in_3_write_data__din),
    .write_data_full_n(mat_C_ch_in_3_write_data__full_n),
    .write_data_write(mat_C_ch_in_3_write_data__write),
    .write_resp_dout(mat_C_ch_in_3_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_3_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_4__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_4___mat_C_ch_in_4__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_4_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_4_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_4_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_4_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_4_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_4_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_4_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_4_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_4_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_4_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_4_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_4_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_4_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_4_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_4_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_4_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_4_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_4_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_4_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_4_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_4_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_4_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_4_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_4_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_4_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_4_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_4_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_4_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_4_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_4_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_4_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_4_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_4_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_4_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_4_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_4_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_4_WVALID),
    .read_addr_din(mat_C_ch_in_4_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_4_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_4_read_addr__write),
    .read_data_dout(mat_C_ch_in_4_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_4_read_data__empty_n),
    .read_data_read(mat_C_ch_in_4_read_data__read),
    .write_addr_din(mat_C_ch_in_4_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_4_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_4_write_addr__write),
    .write_data_din(mat_C_ch_in_4_write_data__din),
    .write_data_full_n(mat_C_ch_in_4_write_data__full_n),
    .write_data_write(mat_C_ch_in_4_write_data__write),
    .write_resp_dout(mat_C_ch_in_4_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_4_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_4_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_5__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_5___mat_C_ch_in_5__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_5_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_5_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_5_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_5_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_5_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_5_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_5_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_5_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_5_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_5_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_5_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_5_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_5_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_5_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_5_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_5_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_5_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_5_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_5_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_5_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_5_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_5_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_5_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_5_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_5_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_5_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_5_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_5_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_5_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_5_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_5_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_5_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_5_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_5_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_5_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_5_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_5_WVALID),
    .read_addr_din(mat_C_ch_in_5_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_5_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_5_read_addr__write),
    .read_data_dout(mat_C_ch_in_5_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_5_read_data__empty_n),
    .read_data_read(mat_C_ch_in_5_read_data__read),
    .write_addr_din(mat_C_ch_in_5_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_5_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_5_write_addr__write),
    .write_data_din(mat_C_ch_in_5_write_data__din),
    .write_data_full_n(mat_C_ch_in_5_write_data__full_n),
    .write_data_write(mat_C_ch_in_5_write_data__write),
    .write_resp_dout(mat_C_ch_in_5_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_5_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_5_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_6__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_6___mat_C_ch_in_6__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_6_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_6_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_6_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_6_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_6_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_6_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_6_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_6_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_6_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_6_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_6_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_6_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_6_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_6_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_6_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_6_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_6_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_6_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_6_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_6_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_6_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_6_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_6_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_6_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_6_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_6_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_6_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_6_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_6_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_6_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_6_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_6_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_6_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_6_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_6_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_6_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_6_WVALID),
    .read_addr_din(mat_C_ch_in_6_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_6_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_6_read_addr__write),
    .read_data_dout(mat_C_ch_in_6_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_6_read_data__empty_n),
    .read_data_read(mat_C_ch_in_6_read_data__read),
    .write_addr_din(mat_C_ch_in_6_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_6_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_6_write_addr__write),
    .write_data_din(mat_C_ch_in_6_write_data__din),
    .write_data_full_n(mat_C_ch_in_6_write_data__full_n),
    .write_data_write(mat_C_ch_in_6_write_data__write),
    .write_resp_dout(mat_C_ch_in_6_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_6_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_6_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_in_7__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_C_7___mat_C_ch_in_7__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_in_7_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_in_7_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_in_7_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_in_7_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_in_7_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_in_7_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_in_7_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_in_7_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_in_7_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_in_7_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_in_7_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_in_7_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_in_7_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_in_7_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_in_7_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_in_7_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_in_7_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_in_7_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_in_7_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_in_7_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_in_7_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_in_7_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_in_7_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_in_7_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_in_7_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_in_7_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_in_7_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_in_7_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_in_7_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_in_7_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_in_7_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_in_7_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_in_7_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_in_7_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_in_7_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_in_7_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_in_7_WVALID),
    .read_addr_din(mat_C_ch_in_7_read_addr__din),
    .read_addr_full_n(mat_C_ch_in_7_read_addr__full_n),
    .read_addr_write(mat_C_ch_in_7_read_addr__write),
    .read_data_dout(mat_C_ch_in_7_read_data__dout),
    .read_data_empty_n(mat_C_ch_in_7_read_data__empty_n),
    .read_data_read(mat_C_ch_in_7_read_data__read),
    .write_addr_din(mat_C_ch_in_7_write_addr__din),
    .write_addr_full_n(mat_C_ch_in_7_write_addr__full_n),
    .write_addr_write(mat_C_ch_in_7_write_addr__write),
    .write_data_din(mat_C_ch_in_7_write_data__din),
    .write_data_full_n(mat_C_ch_in_7_write_data__full_n),
    .write_data_write(mat_C_ch_in_7_write_data__write),
    .write_resp_dout(mat_C_ch_in_7_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_in_7_write_resp__empty_n),
    .write_resp_read(mat_C_ch_in_7_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(32),
    .DataWidthBytesLog(2),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(255)
  )
  edge_list_ptr__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(read_edge_list_ptr_0___edge_list_ptr__q0),
    .m_axi_ARADDR(m_axi_edge_list_ptr_ARADDR),
    .m_axi_ARBURST(m_axi_edge_list_ptr_ARBURST),
    .m_axi_ARCACHE(m_axi_edge_list_ptr_ARCACHE),
    .m_axi_ARID(m_axi_edge_list_ptr_ARID),
    .m_axi_ARLEN(m_axi_edge_list_ptr_ARLEN),
    .m_axi_ARLOCK(m_axi_edge_list_ptr_ARLOCK),
    .m_axi_ARPROT(m_axi_edge_list_ptr_ARPROT),
    .m_axi_ARQOS(m_axi_edge_list_ptr_ARQOS),
    .m_axi_ARREADY(m_axi_edge_list_ptr_ARREADY),
    .m_axi_ARSIZE(m_axi_edge_list_ptr_ARSIZE),
    .m_axi_ARVALID(m_axi_edge_list_ptr_ARVALID),
    .m_axi_AWADDR(m_axi_edge_list_ptr_AWADDR),
    .m_axi_AWBURST(m_axi_edge_list_ptr_AWBURST),
    .m_axi_AWCACHE(m_axi_edge_list_ptr_AWCACHE),
    .m_axi_AWID(m_axi_edge_list_ptr_AWID),
    .m_axi_AWLEN(m_axi_edge_list_ptr_AWLEN),
    .m_axi_AWLOCK(m_axi_edge_list_ptr_AWLOCK),
    .m_axi_AWPROT(m_axi_edge_list_ptr_AWPROT),
    .m_axi_AWQOS(m_axi_edge_list_ptr_AWQOS),
    .m_axi_AWREADY(m_axi_edge_list_ptr_AWREADY),
    .m_axi_AWSIZE(m_axi_edge_list_ptr_AWSIZE),
    .m_axi_AWVALID(m_axi_edge_list_ptr_AWVALID),
    .m_axi_BID(m_axi_edge_list_ptr_BID),
    .m_axi_BREADY(m_axi_edge_list_ptr_BREADY),
    .m_axi_BRESP(m_axi_edge_list_ptr_BRESP),
    .m_axi_BVALID(m_axi_edge_list_ptr_BVALID),
    .m_axi_RDATA(m_axi_edge_list_ptr_RDATA),
    .m_axi_RID(m_axi_edge_list_ptr_RID),
    .m_axi_RLAST(m_axi_edge_list_ptr_RLAST),
    .m_axi_RREADY(m_axi_edge_list_ptr_RREADY),
    .m_axi_RRESP(m_axi_edge_list_ptr_RRESP),
    .m_axi_RVALID(m_axi_edge_list_ptr_RVALID),
    .m_axi_WDATA(m_axi_edge_list_ptr_WDATA),
    .m_axi_WLAST(m_axi_edge_list_ptr_WLAST),
    .m_axi_WREADY(m_axi_edge_list_ptr_WREADY),
    .m_axi_WSTRB(m_axi_edge_list_ptr_WSTRB),
    .m_axi_WVALID(m_axi_edge_list_ptr_WVALID),
    .read_addr_din(edge_list_ptr_read_addr__din),
    .read_addr_full_n(edge_list_ptr_read_addr__full_n),
    .read_addr_write(edge_list_ptr_read_addr__write),
    .read_data_dout(edge_list_ptr_read_data__dout),
    .read_data_empty_n(edge_list_ptr_read_data__empty_n),
    .read_data_read(edge_list_ptr_read_data__read),
    .write_addr_din(edge_list_ptr_write_addr__din),
    .write_addr_full_n(edge_list_ptr_write_addr__full_n),
    .write_addr_write(edge_list_ptr_write_addr__write),
    .write_data_din(edge_list_ptr_write_data__din),
    .write_data_full_n(edge_list_ptr_write_data__full_n),
    .write_data_write(edge_list_ptr_write_data__write),
    .write_resp_dout(edge_list_ptr_write_resp__dout),
    .write_resp_empty_n(edge_list_ptr_write_resp__empty_n),
    .write_resp_read(edge_list_ptr_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_0___mat_C_ch_0__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_0_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_0_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_0_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_0_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_0_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_0_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_0_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_0_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_0_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_0_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_0_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_0_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_0_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_0_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_0_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_0_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_0_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_0_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_0_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_0_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_0_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_0_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_0_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_0_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_0_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_0_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_0_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_0_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_0_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_0_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_0_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_0_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_0_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_0_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_0_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_0_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_0_WVALID),
    .read_addr_din(mat_C_ch_0_read_addr__din),
    .read_addr_full_n(mat_C_ch_0_read_addr__full_n),
    .read_addr_write(mat_C_ch_0_read_addr__write),
    .read_data_dout(mat_C_ch_0_read_data__dout),
    .read_data_empty_n(mat_C_ch_0_read_data__empty_n),
    .read_data_read(mat_C_ch_0_read_data__read),
    .write_addr_din(mat_C_ch_0_write_addr__din),
    .write_addr_full_n(mat_C_ch_0_write_addr__full_n),
    .write_addr_write(mat_C_ch_0_write_addr__write),
    .write_data_din(mat_C_ch_0_write_data__din),
    .write_data_full_n(mat_C_ch_0_write_data__full_n),
    .write_data_write(mat_C_ch_0_write_data__write),
    .write_resp_dout(mat_C_ch_0_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_0_write_resp__empty_n),
    .write_resp_read(mat_C_ch_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_1___mat_C_ch_1__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_1_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_1_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_1_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_1_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_1_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_1_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_1_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_1_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_1_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_1_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_1_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_1_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_1_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_1_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_1_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_1_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_1_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_1_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_1_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_1_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_1_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_1_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_1_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_1_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_1_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_1_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_1_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_1_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_1_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_1_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_1_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_1_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_1_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_1_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_1_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_1_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_1_WVALID),
    .read_addr_din(mat_C_ch_1_read_addr__din),
    .read_addr_full_n(mat_C_ch_1_read_addr__full_n),
    .read_addr_write(mat_C_ch_1_read_addr__write),
    .read_data_dout(mat_C_ch_1_read_data__dout),
    .read_data_empty_n(mat_C_ch_1_read_data__empty_n),
    .read_data_read(mat_C_ch_1_read_data__read),
    .write_addr_din(mat_C_ch_1_write_addr__din),
    .write_addr_full_n(mat_C_ch_1_write_addr__full_n),
    .write_addr_write(mat_C_ch_1_write_addr__write),
    .write_data_din(mat_C_ch_1_write_data__din),
    .write_data_full_n(mat_C_ch_1_write_data__full_n),
    .write_data_write(mat_C_ch_1_write_data__write),
    .write_resp_dout(mat_C_ch_1_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_1_write_resp__empty_n),
    .write_resp_read(mat_C_ch_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_2___mat_C_ch_2__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_2_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_2_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_2_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_2_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_2_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_2_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_2_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_2_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_2_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_2_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_2_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_2_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_2_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_2_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_2_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_2_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_2_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_2_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_2_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_2_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_2_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_2_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_2_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_2_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_2_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_2_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_2_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_2_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_2_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_2_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_2_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_2_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_2_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_2_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_2_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_2_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_2_WVALID),
    .read_addr_din(mat_C_ch_2_read_addr__din),
    .read_addr_full_n(mat_C_ch_2_read_addr__full_n),
    .read_addr_write(mat_C_ch_2_read_addr__write),
    .read_data_dout(mat_C_ch_2_read_data__dout),
    .read_data_empty_n(mat_C_ch_2_read_data__empty_n),
    .read_data_read(mat_C_ch_2_read_data__read),
    .write_addr_din(mat_C_ch_2_write_addr__din),
    .write_addr_full_n(mat_C_ch_2_write_addr__full_n),
    .write_addr_write(mat_C_ch_2_write_addr__write),
    .write_data_din(mat_C_ch_2_write_data__din),
    .write_data_full_n(mat_C_ch_2_write_data__full_n),
    .write_data_write(mat_C_ch_2_write_data__write),
    .write_resp_dout(mat_C_ch_2_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_2_write_resp__empty_n),
    .write_resp_read(mat_C_ch_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_3___mat_C_ch_3__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_3_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_3_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_3_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_3_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_3_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_3_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_3_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_3_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_3_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_3_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_3_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_3_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_3_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_3_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_3_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_3_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_3_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_3_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_3_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_3_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_3_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_3_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_3_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_3_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_3_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_3_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_3_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_3_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_3_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_3_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_3_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_3_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_3_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_3_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_3_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_3_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_3_WVALID),
    .read_addr_din(mat_C_ch_3_read_addr__din),
    .read_addr_full_n(mat_C_ch_3_read_addr__full_n),
    .read_addr_write(mat_C_ch_3_read_addr__write),
    .read_data_dout(mat_C_ch_3_read_data__dout),
    .read_data_empty_n(mat_C_ch_3_read_data__empty_n),
    .read_data_read(mat_C_ch_3_read_data__read),
    .write_addr_din(mat_C_ch_3_write_addr__din),
    .write_addr_full_n(mat_C_ch_3_write_addr__full_n),
    .write_addr_write(mat_C_ch_3_write_addr__write),
    .write_data_din(mat_C_ch_3_write_data__din),
    .write_data_full_n(mat_C_ch_3_write_data__full_n),
    .write_data_write(mat_C_ch_3_write_data__write),
    .write_resp_dout(mat_C_ch_3_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_3_write_resp__empty_n),
    .write_resp_read(mat_C_ch_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_4__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_4___mat_C_ch_4__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_4_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_4_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_4_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_4_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_4_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_4_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_4_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_4_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_4_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_4_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_4_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_4_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_4_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_4_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_4_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_4_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_4_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_4_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_4_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_4_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_4_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_4_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_4_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_4_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_4_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_4_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_4_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_4_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_4_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_4_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_4_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_4_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_4_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_4_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_4_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_4_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_4_WVALID),
    .read_addr_din(mat_C_ch_4_read_addr__din),
    .read_addr_full_n(mat_C_ch_4_read_addr__full_n),
    .read_addr_write(mat_C_ch_4_read_addr__write),
    .read_data_dout(mat_C_ch_4_read_data__dout),
    .read_data_empty_n(mat_C_ch_4_read_data__empty_n),
    .read_data_read(mat_C_ch_4_read_data__read),
    .write_addr_din(mat_C_ch_4_write_addr__din),
    .write_addr_full_n(mat_C_ch_4_write_addr__full_n),
    .write_addr_write(mat_C_ch_4_write_addr__write),
    .write_data_din(mat_C_ch_4_write_data__din),
    .write_data_full_n(mat_C_ch_4_write_data__full_n),
    .write_data_write(mat_C_ch_4_write_data__write),
    .write_resp_dout(mat_C_ch_4_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_4_write_resp__empty_n),
    .write_resp_read(mat_C_ch_4_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_5__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_5___mat_C_ch_5__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_5_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_5_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_5_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_5_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_5_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_5_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_5_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_5_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_5_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_5_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_5_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_5_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_5_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_5_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_5_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_5_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_5_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_5_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_5_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_5_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_5_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_5_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_5_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_5_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_5_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_5_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_5_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_5_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_5_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_5_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_5_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_5_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_5_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_5_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_5_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_5_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_5_WVALID),
    .read_addr_din(mat_C_ch_5_read_addr__din),
    .read_addr_full_n(mat_C_ch_5_read_addr__full_n),
    .read_addr_write(mat_C_ch_5_read_addr__write),
    .read_data_dout(mat_C_ch_5_read_data__dout),
    .read_data_empty_n(mat_C_ch_5_read_data__empty_n),
    .read_data_read(mat_C_ch_5_read_data__read),
    .write_addr_din(mat_C_ch_5_write_addr__din),
    .write_addr_full_n(mat_C_ch_5_write_addr__full_n),
    .write_addr_write(mat_C_ch_5_write_addr__write),
    .write_data_din(mat_C_ch_5_write_data__din),
    .write_data_full_n(mat_C_ch_5_write_data__full_n),
    .write_data_write(mat_C_ch_5_write_data__write),
    .write_resp_dout(mat_C_ch_5_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_5_write_resp__empty_n),
    .write_resp_read(mat_C_ch_5_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_6__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_6___mat_C_ch_6__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_6_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_6_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_6_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_6_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_6_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_6_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_6_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_6_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_6_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_6_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_6_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_6_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_6_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_6_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_6_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_6_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_6_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_6_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_6_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_6_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_6_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_6_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_6_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_6_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_6_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_6_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_6_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_6_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_6_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_6_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_6_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_6_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_6_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_6_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_6_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_6_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_6_WVALID),
    .read_addr_din(mat_C_ch_6_read_addr__din),
    .read_addr_full_n(mat_C_ch_6_read_addr__full_n),
    .read_addr_write(mat_C_ch_6_read_addr__write),
    .read_data_dout(mat_C_ch_6_read_data__dout),
    .read_data_empty_n(mat_C_ch_6_read_data__empty_n),
    .read_data_read(mat_C_ch_6_read_data__read),
    .write_addr_din(mat_C_ch_6_write_addr__din),
    .write_addr_full_n(mat_C_ch_6_write_addr__full_n),
    .write_addr_write(mat_C_ch_6_write_addr__write),
    .write_data_din(mat_C_ch_6_write_data__din),
    .write_data_full_n(mat_C_ch_6_write_data__full_n),
    .write_data_write(mat_C_ch_6_write_data__write),
    .write_resp_dout(mat_C_ch_6_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_6_write_resp__empty_n),
    .write_resp_read(mat_C_ch_6_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  mat_C_ch_7__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .offset(write_C_7___mat_C_ch_7__q0),
    .m_axi_ARADDR(m_axi_mat_C_ch_7_ARADDR),
    .m_axi_ARBURST(m_axi_mat_C_ch_7_ARBURST),
    .m_axi_ARCACHE(m_axi_mat_C_ch_7_ARCACHE),
    .m_axi_ARID(m_axi_mat_C_ch_7_ARID),
    .m_axi_ARLEN(m_axi_mat_C_ch_7_ARLEN),
    .m_axi_ARLOCK(m_axi_mat_C_ch_7_ARLOCK),
    .m_axi_ARPROT(m_axi_mat_C_ch_7_ARPROT),
    .m_axi_ARQOS(m_axi_mat_C_ch_7_ARQOS),
    .m_axi_ARREADY(m_axi_mat_C_ch_7_ARREADY),
    .m_axi_ARSIZE(m_axi_mat_C_ch_7_ARSIZE),
    .m_axi_ARVALID(m_axi_mat_C_ch_7_ARVALID),
    .m_axi_AWADDR(m_axi_mat_C_ch_7_AWADDR),
    .m_axi_AWBURST(m_axi_mat_C_ch_7_AWBURST),
    .m_axi_AWCACHE(m_axi_mat_C_ch_7_AWCACHE),
    .m_axi_AWID(m_axi_mat_C_ch_7_AWID),
    .m_axi_AWLEN(m_axi_mat_C_ch_7_AWLEN),
    .m_axi_AWLOCK(m_axi_mat_C_ch_7_AWLOCK),
    .m_axi_AWPROT(m_axi_mat_C_ch_7_AWPROT),
    .m_axi_AWQOS(m_axi_mat_C_ch_7_AWQOS),
    .m_axi_AWREADY(m_axi_mat_C_ch_7_AWREADY),
    .m_axi_AWSIZE(m_axi_mat_C_ch_7_AWSIZE),
    .m_axi_AWVALID(m_axi_mat_C_ch_7_AWVALID),
    .m_axi_BID(m_axi_mat_C_ch_7_BID),
    .m_axi_BREADY(m_axi_mat_C_ch_7_BREADY),
    .m_axi_BRESP(m_axi_mat_C_ch_7_BRESP),
    .m_axi_BVALID(m_axi_mat_C_ch_7_BVALID),
    .m_axi_RDATA(m_axi_mat_C_ch_7_RDATA),
    .m_axi_RID(m_axi_mat_C_ch_7_RID),
    .m_axi_RLAST(m_axi_mat_C_ch_7_RLAST),
    .m_axi_RREADY(m_axi_mat_C_ch_7_RREADY),
    .m_axi_RRESP(m_axi_mat_C_ch_7_RRESP),
    .m_axi_RVALID(m_axi_mat_C_ch_7_RVALID),
    .m_axi_WDATA(m_axi_mat_C_ch_7_WDATA),
    .m_axi_WLAST(m_axi_mat_C_ch_7_WLAST),
    .m_axi_WREADY(m_axi_mat_C_ch_7_WREADY),
    .m_axi_WSTRB(m_axi_mat_C_ch_7_WSTRB),
    .m_axi_WVALID(m_axi_mat_C_ch_7_WVALID),
    .read_addr_din(mat_C_ch_7_read_addr__din),
    .read_addr_full_n(mat_C_ch_7_read_addr__full_n),
    .read_addr_write(mat_C_ch_7_read_addr__write),
    .read_data_dout(mat_C_ch_7_read_data__dout),
    .read_data_empty_n(mat_C_ch_7_read_data__empty_n),
    .read_data_read(mat_C_ch_7_read_data__read),
    .write_addr_din(mat_C_ch_7_write_addr__din),
    .write_addr_full_n(mat_C_ch_7_write_addr__full_n),
    .write_addr_write(mat_C_ch_7_write_addr__write),
    .write_data_din(mat_C_ch_7_write_data__din),
    .write_data_full_n(mat_C_ch_7_write_data__full_n),
    .write_data_write(mat_C_ch_7_write_data__write),
    .write_resp_dout(mat_C_ch_7_write_resp__dout),
    .write_resp_empty_n(mat_C_ch_7_write_resp__empty_n),
    .write_resp_read(mat_C_ch_7_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) Sextans_fsm
  __tapa_fsm_unit
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .FloatvAddFloatv_0__ap_start(FloatvAddFloatv_0__ap_start),
    .FloatvAddFloatv_1__ap_start(FloatvAddFloatv_1__ap_start),
    .FloatvAddFloatv_2__ap_start(FloatvAddFloatv_2__ap_start),
    .FloatvAddFloatv_3__ap_start(FloatvAddFloatv_3__ap_start),
    .FloatvAddFloatv_4__ap_start(FloatvAddFloatv_4__ap_start),
    .FloatvAddFloatv_5__ap_start(FloatvAddFloatv_5__ap_start),
    .FloatvAddFloatv_6__ap_start(FloatvAddFloatv_6__ap_start),
    .FloatvAddFloatv_7__ap_start(FloatvAddFloatv_7__ap_start),
    .FloatvMultConst_0__ap_start(FloatvMultConst_0__ap_start),
    .FloatvMultConst_0__ap_ready(FloatvMultConst_0__ap_ready),
    .FloatvMultConst_0__ap_done(FloatvMultConst_0__ap_done),
    .FloatvMultConst_0__ap_idle(FloatvMultConst_0__ap_idle),
    .FloatvMultConst_1__ap_start(FloatvMultConst_1__ap_start),
    .FloatvMultConst_1__ap_ready(FloatvMultConst_1__ap_ready),
    .FloatvMultConst_1__ap_done(FloatvMultConst_1__ap_done),
    .FloatvMultConst_1__ap_idle(FloatvMultConst_1__ap_idle),
    .FloatvMultConst_2__ap_start(FloatvMultConst_2__ap_start),
    .FloatvMultConst_2__ap_ready(FloatvMultConst_2__ap_ready),
    .FloatvMultConst_2__ap_done(FloatvMultConst_2__ap_done),
    .FloatvMultConst_2__ap_idle(FloatvMultConst_2__ap_idle),
    .FloatvMultConst_3__ap_start(FloatvMultConst_3__ap_start),
    .FloatvMultConst_3__ap_ready(FloatvMultConst_3__ap_ready),
    .FloatvMultConst_3__ap_done(FloatvMultConst_3__ap_done),
    .FloatvMultConst_3__ap_idle(FloatvMultConst_3__ap_idle),
    .FloatvMultConst_4__ap_start(FloatvMultConst_4__ap_start),
    .FloatvMultConst_4__ap_ready(FloatvMultConst_4__ap_ready),
    .FloatvMultConst_4__ap_done(FloatvMultConst_4__ap_done),
    .FloatvMultConst_4__ap_idle(FloatvMultConst_4__ap_idle),
    .FloatvMultConst_5__ap_start(FloatvMultConst_5__ap_start),
    .FloatvMultConst_5__ap_ready(FloatvMultConst_5__ap_ready),
    .FloatvMultConst_5__ap_done(FloatvMultConst_5__ap_done),
    .FloatvMultConst_5__ap_idle(FloatvMultConst_5__ap_idle),
    .FloatvMultConst_6__ap_start(FloatvMultConst_6__ap_start),
    .FloatvMultConst_6__ap_ready(FloatvMultConst_6__ap_ready),
    .FloatvMultConst_6__ap_done(FloatvMultConst_6__ap_done),
    .FloatvMultConst_6__ap_idle(FloatvMultConst_6__ap_idle),
    .FloatvMultConst_7__ap_start(FloatvMultConst_7__ap_start),
    .FloatvMultConst_7__ap_ready(FloatvMultConst_7__ap_ready),
    .FloatvMultConst_7__ap_done(FloatvMultConst_7__ap_done),
    .FloatvMultConst_7__ap_idle(FloatvMultConst_7__ap_idle),
    .FloatvMultConst_8__ap_start(FloatvMultConst_8__ap_start),
    .FloatvMultConst_8__ap_ready(FloatvMultConst_8__ap_ready),
    .FloatvMultConst_8__ap_done(FloatvMultConst_8__ap_done),
    .FloatvMultConst_8__ap_idle(FloatvMultConst_8__ap_idle),
    .FloatvMultConst_9__ap_start(FloatvMultConst_9__ap_start),
    .FloatvMultConst_9__ap_ready(FloatvMultConst_9__ap_ready),
    .FloatvMultConst_9__ap_done(FloatvMultConst_9__ap_done),
    .FloatvMultConst_9__ap_idle(FloatvMultConst_9__ap_idle),
    .FloatvMultConst_10__ap_start(FloatvMultConst_10__ap_start),
    .FloatvMultConst_10__ap_ready(FloatvMultConst_10__ap_ready),
    .FloatvMultConst_10__ap_done(FloatvMultConst_10__ap_done),
    .FloatvMultConst_10__ap_idle(FloatvMultConst_10__ap_idle),
    .FloatvMultConst_11__ap_start(FloatvMultConst_11__ap_start),
    .FloatvMultConst_11__ap_ready(FloatvMultConst_11__ap_ready),
    .FloatvMultConst_11__ap_done(FloatvMultConst_11__ap_done),
    .FloatvMultConst_11__ap_idle(FloatvMultConst_11__ap_idle),
    .FloatvMultConst_12__ap_start(FloatvMultConst_12__ap_start),
    .FloatvMultConst_12__ap_ready(FloatvMultConst_12__ap_ready),
    .FloatvMultConst_12__ap_done(FloatvMultConst_12__ap_done),
    .FloatvMultConst_12__ap_idle(FloatvMultConst_12__ap_idle),
    .FloatvMultConst_13__ap_start(FloatvMultConst_13__ap_start),
    .FloatvMultConst_13__ap_ready(FloatvMultConst_13__ap_ready),
    .FloatvMultConst_13__ap_done(FloatvMultConst_13__ap_done),
    .FloatvMultConst_13__ap_idle(FloatvMultConst_13__ap_idle),
    .FloatvMultConst_14__ap_start(FloatvMultConst_14__ap_start),
    .FloatvMultConst_14__ap_ready(FloatvMultConst_14__ap_ready),
    .FloatvMultConst_14__ap_done(FloatvMultConst_14__ap_done),
    .FloatvMultConst_14__ap_idle(FloatvMultConst_14__ap_idle),
    .FloatvMultConst_15__ap_start(FloatvMultConst_15__ap_start),
    .FloatvMultConst_15__ap_ready(FloatvMultConst_15__ap_ready),
    .FloatvMultConst_15__ap_done(FloatvMultConst_15__ap_done),
    .FloatvMultConst_15__ap_idle(FloatvMultConst_15__ap_idle),
    .Merger_0__ap_start(Merger_0__ap_start),
    .Merger_1__ap_start(Merger_1__ap_start),
    .Merger_2__ap_start(Merger_2__ap_start),
    .Merger_3__ap_start(Merger_3__ap_start),
    .Merger_4__ap_start(Merger_4__ap_start),
    .Merger_5__ap_start(Merger_5__ap_start),
    .Merger_6__ap_start(Merger_6__ap_start),
    .Merger_7__ap_start(Merger_7__ap_start),
    .PEG_Bmtx_0__ap_start(PEG_Bmtx_0__ap_start),
    .PEG_Bmtx_0__ap_ready(PEG_Bmtx_0__ap_ready),
    .PEG_Bmtx_0__ap_done(PEG_Bmtx_0__ap_done),
    .PEG_Bmtx_0__ap_idle(PEG_Bmtx_0__ap_idle),
    .PEG_Bmtx_1__ap_start(PEG_Bmtx_1__ap_start),
    .PEG_Bmtx_1__ap_ready(PEG_Bmtx_1__ap_ready),
    .PEG_Bmtx_1__ap_done(PEG_Bmtx_1__ap_done),
    .PEG_Bmtx_1__ap_idle(PEG_Bmtx_1__ap_idle),
    .PEG_Bmtx_2__ap_start(PEG_Bmtx_2__ap_start),
    .PEG_Bmtx_2__ap_ready(PEG_Bmtx_2__ap_ready),
    .PEG_Bmtx_2__ap_done(PEG_Bmtx_2__ap_done),
    .PEG_Bmtx_2__ap_idle(PEG_Bmtx_2__ap_idle),
    .PEG_Bmtx_3__ap_start(PEG_Bmtx_3__ap_start),
    .PEG_Bmtx_3__ap_ready(PEG_Bmtx_3__ap_ready),
    .PEG_Bmtx_3__ap_done(PEG_Bmtx_3__ap_done),
    .PEG_Bmtx_3__ap_idle(PEG_Bmtx_3__ap_idle),
    .PEG_Bmtx_4__ap_start(PEG_Bmtx_4__ap_start),
    .PEG_Bmtx_4__ap_ready(PEG_Bmtx_4__ap_ready),
    .PEG_Bmtx_4__ap_done(PEG_Bmtx_4__ap_done),
    .PEG_Bmtx_4__ap_idle(PEG_Bmtx_4__ap_idle),
    .PEG_Bmtx_5__ap_start(PEG_Bmtx_5__ap_start),
    .PEG_Bmtx_5__ap_ready(PEG_Bmtx_5__ap_ready),
    .PEG_Bmtx_5__ap_done(PEG_Bmtx_5__ap_done),
    .PEG_Bmtx_5__ap_idle(PEG_Bmtx_5__ap_idle),
    .PEG_Bmtx_6__ap_start(PEG_Bmtx_6__ap_start),
    .PEG_Bmtx_6__ap_ready(PEG_Bmtx_6__ap_ready),
    .PEG_Bmtx_6__ap_done(PEG_Bmtx_6__ap_done),
    .PEG_Bmtx_6__ap_idle(PEG_Bmtx_6__ap_idle),
    .PEG_Bmtx_7__ap_start(PEG_Bmtx_7__ap_start),
    .PEG_Bmtx_7__ap_ready(PEG_Bmtx_7__ap_ready),
    .PEG_Bmtx_7__ap_done(PEG_Bmtx_7__ap_done),
    .PEG_Bmtx_7__ap_idle(PEG_Bmtx_7__ap_idle),
    .PEG_Bmtx_8__ap_start(PEG_Bmtx_8__ap_start),
    .PEG_Bmtx_8__ap_ready(PEG_Bmtx_8__ap_ready),
    .PEG_Bmtx_8__ap_done(PEG_Bmtx_8__ap_done),
    .PEG_Bmtx_8__ap_idle(PEG_Bmtx_8__ap_idle),
    .PEG_Bmtx_9__ap_start(PEG_Bmtx_9__ap_start),
    .PEG_Bmtx_9__ap_ready(PEG_Bmtx_9__ap_ready),
    .PEG_Bmtx_9__ap_done(PEG_Bmtx_9__ap_done),
    .PEG_Bmtx_9__ap_idle(PEG_Bmtx_9__ap_idle),
    .PEG_Bmtx_10__ap_start(PEG_Bmtx_10__ap_start),
    .PEG_Bmtx_10__ap_ready(PEG_Bmtx_10__ap_ready),
    .PEG_Bmtx_10__ap_done(PEG_Bmtx_10__ap_done),
    .PEG_Bmtx_10__ap_idle(PEG_Bmtx_10__ap_idle),
    .PEG_Bmtx_11__ap_start(PEG_Bmtx_11__ap_start),
    .PEG_Bmtx_11__ap_ready(PEG_Bmtx_11__ap_ready),
    .PEG_Bmtx_11__ap_done(PEG_Bmtx_11__ap_done),
    .PEG_Bmtx_11__ap_idle(PEG_Bmtx_11__ap_idle),
    .PEG_Bmtx_12__ap_start(PEG_Bmtx_12__ap_start),
    .PEG_Bmtx_12__ap_ready(PEG_Bmtx_12__ap_ready),
    .PEG_Bmtx_12__ap_done(PEG_Bmtx_12__ap_done),
    .PEG_Bmtx_12__ap_idle(PEG_Bmtx_12__ap_idle),
    .PEG_Bmtx_13__ap_start(PEG_Bmtx_13__ap_start),
    .PEG_Bmtx_13__ap_ready(PEG_Bmtx_13__ap_ready),
    .PEG_Bmtx_13__ap_done(PEG_Bmtx_13__ap_done),
    .PEG_Bmtx_13__ap_idle(PEG_Bmtx_13__ap_idle),
    .PEG_Bmtx_14__ap_start(PEG_Bmtx_14__ap_start),
    .PEG_Bmtx_14__ap_ready(PEG_Bmtx_14__ap_ready),
    .PEG_Bmtx_14__ap_done(PEG_Bmtx_14__ap_done),
    .PEG_Bmtx_14__ap_idle(PEG_Bmtx_14__ap_idle),
    .PEG_Bmtx_15__ap_start(PEG_Bmtx_15__ap_start),
    .PEG_Bmtx_15__ap_ready(PEG_Bmtx_15__ap_ready),
    .PEG_Bmtx_15__ap_done(PEG_Bmtx_15__ap_done),
    .PEG_Bmtx_15__ap_idle(PEG_Bmtx_15__ap_idle),
    .PEG_Cmtx_0__ap_start(PEG_Cmtx_0__ap_start),
    .PEG_Cmtx_0__ap_ready(PEG_Cmtx_0__ap_ready),
    .PEG_Cmtx_0__ap_done(PEG_Cmtx_0__ap_done),
    .PEG_Cmtx_0__ap_idle(PEG_Cmtx_0__ap_idle),
    .PEG_Cmtx_1__ap_start(PEG_Cmtx_1__ap_start),
    .PEG_Cmtx_1__ap_ready(PEG_Cmtx_1__ap_ready),
    .PEG_Cmtx_1__ap_done(PEG_Cmtx_1__ap_done),
    .PEG_Cmtx_1__ap_idle(PEG_Cmtx_1__ap_idle),
    .PEG_Cmtx_2__ap_start(PEG_Cmtx_2__ap_start),
    .PEG_Cmtx_2__ap_ready(PEG_Cmtx_2__ap_ready),
    .PEG_Cmtx_2__ap_done(PEG_Cmtx_2__ap_done),
    .PEG_Cmtx_2__ap_idle(PEG_Cmtx_2__ap_idle),
    .PEG_Cmtx_3__ap_start(PEG_Cmtx_3__ap_start),
    .PEG_Cmtx_3__ap_ready(PEG_Cmtx_3__ap_ready),
    .PEG_Cmtx_3__ap_done(PEG_Cmtx_3__ap_done),
    .PEG_Cmtx_3__ap_idle(PEG_Cmtx_3__ap_idle),
    .PEG_Cmtx_4__ap_start(PEG_Cmtx_4__ap_start),
    .PEG_Cmtx_4__ap_ready(PEG_Cmtx_4__ap_ready),
    .PEG_Cmtx_4__ap_done(PEG_Cmtx_4__ap_done),
    .PEG_Cmtx_4__ap_idle(PEG_Cmtx_4__ap_idle),
    .PEG_Cmtx_5__ap_start(PEG_Cmtx_5__ap_start),
    .PEG_Cmtx_5__ap_ready(PEG_Cmtx_5__ap_ready),
    .PEG_Cmtx_5__ap_done(PEG_Cmtx_5__ap_done),
    .PEG_Cmtx_5__ap_idle(PEG_Cmtx_5__ap_idle),
    .PEG_Cmtx_6__ap_start(PEG_Cmtx_6__ap_start),
    .PEG_Cmtx_6__ap_ready(PEG_Cmtx_6__ap_ready),
    .PEG_Cmtx_6__ap_done(PEG_Cmtx_6__ap_done),
    .PEG_Cmtx_6__ap_idle(PEG_Cmtx_6__ap_idle),
    .PEG_Cmtx_7__ap_start(PEG_Cmtx_7__ap_start),
    .PEG_Cmtx_7__ap_ready(PEG_Cmtx_7__ap_ready),
    .PEG_Cmtx_7__ap_done(PEG_Cmtx_7__ap_done),
    .PEG_Cmtx_7__ap_idle(PEG_Cmtx_7__ap_idle),
    .PEG_Cmtx_8__ap_start(PEG_Cmtx_8__ap_start),
    .PEG_Cmtx_8__ap_ready(PEG_Cmtx_8__ap_ready),
    .PEG_Cmtx_8__ap_done(PEG_Cmtx_8__ap_done),
    .PEG_Cmtx_8__ap_idle(PEG_Cmtx_8__ap_idle),
    .PEG_Cmtx_9__ap_start(PEG_Cmtx_9__ap_start),
    .PEG_Cmtx_9__ap_ready(PEG_Cmtx_9__ap_ready),
    .PEG_Cmtx_9__ap_done(PEG_Cmtx_9__ap_done),
    .PEG_Cmtx_9__ap_idle(PEG_Cmtx_9__ap_idle),
    .PEG_Cmtx_10__ap_start(PEG_Cmtx_10__ap_start),
    .PEG_Cmtx_10__ap_ready(PEG_Cmtx_10__ap_ready),
    .PEG_Cmtx_10__ap_done(PEG_Cmtx_10__ap_done),
    .PEG_Cmtx_10__ap_idle(PEG_Cmtx_10__ap_idle),
    .PEG_Cmtx_11__ap_start(PEG_Cmtx_11__ap_start),
    .PEG_Cmtx_11__ap_ready(PEG_Cmtx_11__ap_ready),
    .PEG_Cmtx_11__ap_done(PEG_Cmtx_11__ap_done),
    .PEG_Cmtx_11__ap_idle(PEG_Cmtx_11__ap_idle),
    .PEG_Cmtx_12__ap_start(PEG_Cmtx_12__ap_start),
    .PEG_Cmtx_12__ap_ready(PEG_Cmtx_12__ap_ready),
    .PEG_Cmtx_12__ap_done(PEG_Cmtx_12__ap_done),
    .PEG_Cmtx_12__ap_idle(PEG_Cmtx_12__ap_idle),
    .PEG_Cmtx_13__ap_start(PEG_Cmtx_13__ap_start),
    .PEG_Cmtx_13__ap_ready(PEG_Cmtx_13__ap_ready),
    .PEG_Cmtx_13__ap_done(PEG_Cmtx_13__ap_done),
    .PEG_Cmtx_13__ap_idle(PEG_Cmtx_13__ap_idle),
    .PEG_Cmtx_14__ap_start(PEG_Cmtx_14__ap_start),
    .PEG_Cmtx_14__ap_ready(PEG_Cmtx_14__ap_ready),
    .PEG_Cmtx_14__ap_done(PEG_Cmtx_14__ap_done),
    .PEG_Cmtx_14__ap_idle(PEG_Cmtx_14__ap_idle),
    .PEG_Cmtx_15__ap_start(PEG_Cmtx_15__ap_start),
    .PEG_Cmtx_15__ap_ready(PEG_Cmtx_15__ap_ready),
    .PEG_Cmtx_15__ap_done(PEG_Cmtx_15__ap_done),
    .PEG_Cmtx_15__ap_idle(PEG_Cmtx_15__ap_idle),
    .Scatter_1_2_0__ap_start(Scatter_1_2_0__ap_start),
    .Scatter_1_2_1__ap_start(Scatter_1_2_1__ap_start),
    .Scatter_1_2_2__ap_start(Scatter_1_2_2__ap_start),
    .Scatter_1_2_3__ap_start(Scatter_1_2_3__ap_start),
    .Scatter_1_2_4__ap_start(Scatter_1_2_4__ap_start),
    .Scatter_1_2_5__ap_start(Scatter_1_2_5__ap_start),
    .Scatter_1_2_6__ap_start(Scatter_1_2_6__ap_start),
    .Scatter_1_2_7__ap_start(Scatter_1_2_7__ap_start),
    .black_hole_float_v16_0__ap_start(black_hole_float_v16_0__ap_start),
    .black_hole_float_v16_1__ap_start(black_hole_float_v16_1__ap_start),
    .black_hole_float_v16_2__ap_start(black_hole_float_v16_2__ap_start),
    .black_hole_float_v16_3__ap_start(black_hole_float_v16_3__ap_start),
    .black_hole_int_0__ap_start(black_hole_int_0__ap_start),
    .black_hole_int_1__ap_start(black_hole_int_1__ap_start),
    .read_A_0__ap_start(read_A_0__ap_start),
    .read_A_0__ap_ready(read_A_0__ap_ready),
    .read_A_0__ap_done(read_A_0__ap_done),
    .read_A_0__ap_idle(read_A_0__ap_idle),
    .read_A_1__ap_start(read_A_1__ap_start),
    .read_A_1__ap_ready(read_A_1__ap_ready),
    .read_A_1__ap_done(read_A_1__ap_done),
    .read_A_1__ap_idle(read_A_1__ap_idle),
    .read_A_2__ap_start(read_A_2__ap_start),
    .read_A_2__ap_ready(read_A_2__ap_ready),
    .read_A_2__ap_done(read_A_2__ap_done),
    .read_A_2__ap_idle(read_A_2__ap_idle),
    .read_A_3__ap_start(read_A_3__ap_start),
    .read_A_3__ap_ready(read_A_3__ap_ready),
    .read_A_3__ap_done(read_A_3__ap_done),
    .read_A_3__ap_idle(read_A_3__ap_idle),
    .read_A_4__ap_start(read_A_4__ap_start),
    .read_A_4__ap_ready(read_A_4__ap_ready),
    .read_A_4__ap_done(read_A_4__ap_done),
    .read_A_4__ap_idle(read_A_4__ap_idle),
    .read_A_5__ap_start(read_A_5__ap_start),
    .read_A_5__ap_ready(read_A_5__ap_ready),
    .read_A_5__ap_done(read_A_5__ap_done),
    .read_A_5__ap_idle(read_A_5__ap_idle),
    .read_A_6__ap_start(read_A_6__ap_start),
    .read_A_6__ap_ready(read_A_6__ap_ready),
    .read_A_6__ap_done(read_A_6__ap_done),
    .read_A_6__ap_idle(read_A_6__ap_idle),
    .read_A_7__ap_start(read_A_7__ap_start),
    .read_A_7__ap_ready(read_A_7__ap_ready),
    .read_A_7__ap_done(read_A_7__ap_done),
    .read_A_7__ap_idle(read_A_7__ap_idle),
    .read_B_0__ap_start(read_B_0__ap_start),
    .read_B_0__ap_ready(read_B_0__ap_ready),
    .read_B_0__ap_done(read_B_0__ap_done),
    .read_B_0__ap_idle(read_B_0__ap_idle),
    .read_B_1__ap_start(read_B_1__ap_start),
    .read_B_1__ap_ready(read_B_1__ap_ready),
    .read_B_1__ap_done(read_B_1__ap_done),
    .read_B_1__ap_idle(read_B_1__ap_idle),
    .read_B_2__ap_start(read_B_2__ap_start),
    .read_B_2__ap_ready(read_B_2__ap_ready),
    .read_B_2__ap_done(read_B_2__ap_done),
    .read_B_2__ap_idle(read_B_2__ap_idle),
    .read_B_3__ap_start(read_B_3__ap_start),
    .read_B_3__ap_ready(read_B_3__ap_ready),
    .read_B_3__ap_done(read_B_3__ap_done),
    .read_B_3__ap_idle(read_B_3__ap_idle),
    .read_C_0__ap_start(read_C_0__ap_start),
    .read_C_0__ap_ready(read_C_0__ap_ready),
    .read_C_0__ap_done(read_C_0__ap_done),
    .read_C_0__ap_idle(read_C_0__ap_idle),
    .read_C_1__ap_start(read_C_1__ap_start),
    .read_C_1__ap_ready(read_C_1__ap_ready),
    .read_C_1__ap_done(read_C_1__ap_done),
    .read_C_1__ap_idle(read_C_1__ap_idle),
    .read_C_2__ap_start(read_C_2__ap_start),
    .read_C_2__ap_ready(read_C_2__ap_ready),
    .read_C_2__ap_done(read_C_2__ap_done),
    .read_C_2__ap_idle(read_C_2__ap_idle),
    .read_C_3__ap_start(read_C_3__ap_start),
    .read_C_3__ap_ready(read_C_3__ap_ready),
    .read_C_3__ap_done(read_C_3__ap_done),
    .read_C_3__ap_idle(read_C_3__ap_idle),
    .read_C_4__ap_start(read_C_4__ap_start),
    .read_C_4__ap_ready(read_C_4__ap_ready),
    .read_C_4__ap_done(read_C_4__ap_done),
    .read_C_4__ap_idle(read_C_4__ap_idle),
    .read_C_5__ap_start(read_C_5__ap_start),
    .read_C_5__ap_ready(read_C_5__ap_ready),
    .read_C_5__ap_done(read_C_5__ap_done),
    .read_C_5__ap_idle(read_C_5__ap_idle),
    .read_C_6__ap_start(read_C_6__ap_start),
    .read_C_6__ap_ready(read_C_6__ap_ready),
    .read_C_6__ap_done(read_C_6__ap_done),
    .read_C_6__ap_idle(read_C_6__ap_idle),
    .read_C_7__ap_start(read_C_7__ap_start),
    .read_C_7__ap_ready(read_C_7__ap_ready),
    .read_C_7__ap_done(read_C_7__ap_done),
    .read_C_7__ap_idle(read_C_7__ap_idle),
    .read_edge_list_ptr_0__ap_start(read_edge_list_ptr_0__ap_start),
    .read_edge_list_ptr_0__ap_ready(read_edge_list_ptr_0__ap_ready),
    .read_edge_list_ptr_0__ap_done(read_edge_list_ptr_0__ap_done),
    .read_edge_list_ptr_0__ap_idle(read_edge_list_ptr_0__ap_idle),
    .write_C_0__ap_start(write_C_0__ap_start),
    .write_C_0__ap_ready(write_C_0__ap_ready),
    .write_C_0__ap_done(write_C_0__ap_done),
    .write_C_0__ap_idle(write_C_0__ap_idle),
    .write_C_1__ap_start(write_C_1__ap_start),
    .write_C_1__ap_ready(write_C_1__ap_ready),
    .write_C_1__ap_done(write_C_1__ap_done),
    .write_C_1__ap_idle(write_C_1__ap_idle),
    .write_C_2__ap_start(write_C_2__ap_start),
    .write_C_2__ap_ready(write_C_2__ap_ready),
    .write_C_2__ap_done(write_C_2__ap_done),
    .write_C_2__ap_idle(write_C_2__ap_idle),
    .write_C_3__ap_start(write_C_3__ap_start),
    .write_C_3__ap_ready(write_C_3__ap_ready),
    .write_C_3__ap_done(write_C_3__ap_done),
    .write_C_3__ap_idle(write_C_3__ap_idle),
    .write_C_4__ap_start(write_C_4__ap_start),
    .write_C_4__ap_ready(write_C_4__ap_ready),
    .write_C_4__ap_done(write_C_4__ap_done),
    .write_C_4__ap_idle(write_C_4__ap_idle),
    .write_C_5__ap_start(write_C_5__ap_start),
    .write_C_5__ap_ready(write_C_5__ap_ready),
    .write_C_5__ap_done(write_C_5__ap_done),
    .write_C_5__ap_idle(write_C_5__ap_idle),
    .write_C_6__ap_start(write_C_6__ap_start),
    .write_C_6__ap_ready(write_C_6__ap_ready),
    .write_C_6__ap_done(write_C_6__ap_done),
    .write_C_6__ap_idle(write_C_6__ap_idle),
    .write_C_7__ap_start(write_C_7__ap_start),
    .write_C_7__ap_ready(write_C_7__ap_ready),
    .write_C_7__ap_done(write_C_7__ap_done),
    .write_C_7__ap_idle(write_C_7__ap_idle)
  );

  assign ap_rst_n_inv = (~ap_rst_n);
  assign FloatvMultConst_0___M__q0 = M;
  assign FloatvMultConst_0___P_N__q0 = P_N;
  assign FloatvMultConst_0___beta_u__q0 = beta_u;
  assign FloatvMultConst_1___M__q0 = M;
  assign FloatvMultConst_1___P_N__q0 = P_N;
  assign FloatvMultConst_1___beta_u__q0 = beta_u;
  assign FloatvMultConst_2___M__q0 = M;
  assign FloatvMultConst_2___P_N__q0 = P_N;
  assign FloatvMultConst_2___beta_u__q0 = beta_u;
  assign FloatvMultConst_3___M__q0 = M;
  assign FloatvMultConst_3___P_N__q0 = P_N;
  assign FloatvMultConst_3___beta_u__q0 = beta_u;
  assign FloatvMultConst_4___M__q0 = M;
  assign FloatvMultConst_4___P_N__q0 = P_N;
  assign FloatvMultConst_4___beta_u__q0 = beta_u;
  assign FloatvMultConst_5___M__q0 = M;
  assign FloatvMultConst_5___P_N__q0 = P_N;
  assign FloatvMultConst_5___beta_u__q0 = beta_u;
  assign FloatvMultConst_6___M__q0 = M;
  assign FloatvMultConst_6___P_N__q0 = P_N;
  assign FloatvMultConst_6___beta_u__q0 = beta_u;
  assign FloatvMultConst_7___M__q0 = M;
  assign FloatvMultConst_7___P_N__q0 = P_N;
  assign FloatvMultConst_7___beta_u__q0 = beta_u;
  assign FloatvMultConst_8___M__q0 = M;
  assign FloatvMultConst_8___P_N__q0 = P_N;
  assign FloatvMultConst_8___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_9___M__q0 = M;
  assign FloatvMultConst_9___P_N__q0 = P_N;
  assign FloatvMultConst_9___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_10___M__q0 = M;
  assign FloatvMultConst_10___P_N__q0 = P_N;
  assign FloatvMultConst_10___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_11___M__q0 = M;
  assign FloatvMultConst_11___P_N__q0 = P_N;
  assign FloatvMultConst_11___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_12___M__q0 = M;
  assign FloatvMultConst_12___P_N__q0 = P_N;
  assign FloatvMultConst_12___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_13___M__q0 = M;
  assign FloatvMultConst_13___P_N__q0 = P_N;
  assign FloatvMultConst_13___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_14___M__q0 = M;
  assign FloatvMultConst_14___P_N__q0 = P_N;
  assign FloatvMultConst_14___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_15___M__q0 = M;
  assign FloatvMultConst_15___P_N__q0 = P_N;
  assign FloatvMultConst_15___alpha_u__q0 = alpha_u;
  assign read_A_0___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_0___P_N__q0 = P_N;
  assign read_A_0___edge_list_ch_0__q0 = edge_list_ch_0;
  assign read_A_1___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_1___P_N__q0 = P_N;
  assign read_A_1___edge_list_ch_1__q0 = edge_list_ch_1;
  assign read_A_2___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_2___P_N__q0 = P_N;
  assign read_A_2___edge_list_ch_2__q0 = edge_list_ch_2;
  assign read_A_3___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_3___P_N__q0 = P_N;
  assign read_A_3___edge_list_ch_3__q0 = edge_list_ch_3;
  assign read_A_4___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_4___P_N__q0 = P_N;
  assign read_A_4___edge_list_ch_4__q0 = edge_list_ch_4;
  assign read_A_5___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_5___P_N__q0 = P_N;
  assign read_A_5___edge_list_ch_5__q0 = edge_list_ch_5;
  assign read_A_6___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_6___P_N__q0 = P_N;
  assign read_A_6___edge_list_ch_6__q0 = edge_list_ch_6;
  assign read_A_7___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_7___P_N__q0 = P_N;
  assign read_A_7___edge_list_ch_7__q0 = edge_list_ch_7;
  assign read_B_0___K__q0 = K;
  assign read_B_0___P_N__q0 = P_N;
  assign read_B_0___mat_B_ch_0__q0 = mat_B_ch_0;
  assign read_B_1___K__q0 = K;
  assign read_B_1___P_N__q0 = P_N;
  assign read_B_1___mat_B_ch_1__q0 = mat_B_ch_1;
  assign read_B_2___K__q0 = K;
  assign read_B_2___P_N__q0 = P_N;
  assign read_B_2___mat_B_ch_2__q0 = mat_B_ch_2;
  assign read_B_3___K__q0 = K;
  assign read_B_3___P_N__q0 = P_N;
  assign read_B_3___mat_B_ch_3__q0 = mat_B_ch_3;
  assign read_C_0___M__q0 = M;
  assign read_C_0___P_N__q0 = P_N;
  assign read_C_0___mat_C_ch_in_0__q0 = mat_C_ch_in_0;
  assign read_C_1___M__q0 = M;
  assign read_C_1___P_N__q0 = P_N;
  assign read_C_1___mat_C_ch_in_1__q0 = mat_C_ch_in_1;
  assign read_C_2___M__q0 = M;
  assign read_C_2___P_N__q0 = P_N;
  assign read_C_2___mat_C_ch_in_2__q0 = mat_C_ch_in_2;
  assign read_C_3___M__q0 = M;
  assign read_C_3___P_N__q0 = P_N;
  assign read_C_3___mat_C_ch_in_3__q0 = mat_C_ch_in_3;
  assign read_C_4___M__q0 = M;
  assign read_C_4___P_N__q0 = P_N;
  assign read_C_4___mat_C_ch_in_4__q0 = mat_C_ch_in_4;
  assign read_C_5___M__q0 = M;
  assign read_C_5___P_N__q0 = P_N;
  assign read_C_5___mat_C_ch_in_5__q0 = mat_C_ch_in_5;
  assign read_C_6___M__q0 = M;
  assign read_C_6___P_N__q0 = P_N;
  assign read_C_6___mat_C_ch_in_6__q0 = mat_C_ch_in_6;
  assign read_C_7___M__q0 = M;
  assign read_C_7___P_N__q0 = P_N;
  assign read_C_7___mat_C_ch_in_7__q0 = mat_C_ch_in_7;
  assign read_edge_list_ptr_0___K__q0 = K;
  assign read_edge_list_ptr_0___M__q0 = M;
  assign read_edge_list_ptr_0___NUM_ITE__q0 = NUM_ITE;
  assign read_edge_list_ptr_0___P_N__q0 = P_N;
  assign read_edge_list_ptr_0___edge_list_ptr__q0 = edge_list_ptr;
  assign write_C_0___mat_C_ch_0__q0 = mat_C_ch_0;
  assign write_C_1___mat_C_ch_1__q0 = mat_C_ch_1;
  assign write_C_2___mat_C_ch_2__q0 = mat_C_ch_2;
  assign write_C_3___mat_C_ch_3__q0 = mat_C_ch_3;
  assign write_C_4___mat_C_ch_4__q0 = mat_C_ch_4;
  assign write_C_5___mat_C_ch_5__q0 = mat_C_ch_5;
  assign write_C_6___mat_C_ch_6__q0 = mat_C_ch_6;
  assign write_C_7___mat_C_ch_7__q0 = mat_C_ch_7;

endmodule
