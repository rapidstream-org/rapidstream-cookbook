

module unikernel_fsm
(
  ap_clk,
  ap_rst_n,
  ap_start,
  ap_ready,
  ap_done,
  ap_idle,
  SEIDEL2D_0__ap_start,
  SEIDEL2D_0__ap_ready,
  SEIDEL2D_0__ap_done,
  SEIDEL2D_0__ap_idle,
  SEIDEL2D_1__ap_start,
  SEIDEL2D_1__ap_ready,
  SEIDEL2D_1__ap_done,
  SEIDEL2D_1__ap_idle,
  SEIDEL2D_2__ap_start,
  SEIDEL2D_2__ap_ready,
  SEIDEL2D_2__ap_done,
  SEIDEL2D_2__ap_idle,
  SEIDEL2D_3__ap_start,
  SEIDEL2D_3__ap_ready,
  SEIDEL2D_3__ap_done,
  SEIDEL2D_3__ap_idle,
  SEIDEL2D_4__ap_start,
  SEIDEL2D_4__ap_ready,
  SEIDEL2D_4__ap_done,
  SEIDEL2D_4__ap_idle,
  SEIDEL2D_5__ap_start,
  SEIDEL2D_5__ap_ready,
  SEIDEL2D_5__ap_done,
  SEIDEL2D_5__ap_idle,
  SEIDEL2D_6__ap_start,
  SEIDEL2D_6__ap_ready,
  SEIDEL2D_6__ap_done,
  SEIDEL2D_6__ap_idle,
  SEIDEL2D_7__ap_start,
  SEIDEL2D_7__ap_ready,
  SEIDEL2D_7__ap_done,
  SEIDEL2D_7__ap_idle,
  SEIDEL2D_8__ap_start,
  SEIDEL2D_8__ap_ready,
  SEIDEL2D_8__ap_done,
  SEIDEL2D_8__ap_idle,
  SEIDEL2D_9__ap_start,
  SEIDEL2D_9__ap_ready,
  SEIDEL2D_9__ap_done,
  SEIDEL2D_9__ap_idle,
  SEIDEL2D_10__ap_start,
  SEIDEL2D_10__ap_ready,
  SEIDEL2D_10__ap_done,
  SEIDEL2D_10__ap_idle,
  SEIDEL2D_11__ap_start,
  SEIDEL2D_11__ap_ready,
  SEIDEL2D_11__ap_done,
  SEIDEL2D_11__ap_idle,
  inter_kernel_0__ap_start,
  inter_kernel_0__ap_ready,
  inter_kernel_0__ap_done,
  inter_kernel_0__ap_idle,
  inter_kernel_1__ap_start,
  inter_kernel_1__ap_ready,
  inter_kernel_1__ap_done,
  inter_kernel_1__ap_idle,
  inter_kernel_2__ap_start,
  inter_kernel_2__ap_ready,
  inter_kernel_2__ap_done,
  inter_kernel_2__ap_idle,
  inter_kernel_3__ap_start,
  inter_kernel_3__ap_ready,
  inter_kernel_3__ap_done,
  inter_kernel_3__ap_idle,
  inter_kernel_4__ap_start,
  inter_kernel_4__ap_ready,
  inter_kernel_4__ap_done,
  inter_kernel_4__ap_idle,
  inter_kernel_5__ap_start,
  inter_kernel_5__ap_ready,
  inter_kernel_5__ap_done,
  inter_kernel_5__ap_idle,
  inter_kernel_6__ap_start,
  inter_kernel_6__ap_ready,
  inter_kernel_6__ap_done,
  inter_kernel_6__ap_idle,
  inter_kernel_7__ap_start,
  inter_kernel_7__ap_ready,
  inter_kernel_7__ap_done,
  inter_kernel_7__ap_idle,
  inter_kernel_8__ap_start,
  inter_kernel_8__ap_ready,
  inter_kernel_8__ap_done,
  inter_kernel_8__ap_idle,
  inter_kernel_9__ap_start,
  inter_kernel_9__ap_ready,
  inter_kernel_9__ap_done,
  inter_kernel_9__ap_idle,
  inter_kernel_10__ap_start,
  inter_kernel_10__ap_ready,
  inter_kernel_10__ap_done,
  inter_kernel_10__ap_idle,
  inter_kernel_11__ap_start,
  inter_kernel_11__ap_ready,
  inter_kernel_11__ap_done,
  inter_kernel_11__ap_idle
);

  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_AP_CTRL = "unikernel.ap_start" *)input ap_start;
  (* RS_AP_CTRL = "unikernel.ap_ready" *)output ap_ready;
  (* RS_FF = "unikernel__ap_done" *)output ap_done;
  (* RS_FF = "unikernel__ap_idle" *)output ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_0.ap_start" *)output SEIDEL2D_0__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_0.ap_ready" *)input SEIDEL2D_0__ap_ready;
  (* RS_FF = "SEIDEL2D_0__ap_done" *)input SEIDEL2D_0__ap_done;
  (* RS_FF = "SEIDEL2D_0__ap_idle" *)input SEIDEL2D_0__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_1.ap_start" *)output SEIDEL2D_1__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_1.ap_ready" *)input SEIDEL2D_1__ap_ready;
  (* RS_FF = "SEIDEL2D_1__ap_done" *)input SEIDEL2D_1__ap_done;
  (* RS_FF = "SEIDEL2D_1__ap_idle" *)input SEIDEL2D_1__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_2.ap_start" *)output SEIDEL2D_2__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_2.ap_ready" *)input SEIDEL2D_2__ap_ready;
  (* RS_FF = "SEIDEL2D_2__ap_done" *)input SEIDEL2D_2__ap_done;
  (* RS_FF = "SEIDEL2D_2__ap_idle" *)input SEIDEL2D_2__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_3.ap_start" *)output SEIDEL2D_3__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_3.ap_ready" *)input SEIDEL2D_3__ap_ready;
  (* RS_FF = "SEIDEL2D_3__ap_done" *)input SEIDEL2D_3__ap_done;
  (* RS_FF = "SEIDEL2D_3__ap_idle" *)input SEIDEL2D_3__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_4.ap_start" *)output SEIDEL2D_4__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_4.ap_ready" *)input SEIDEL2D_4__ap_ready;
  (* RS_FF = "SEIDEL2D_4__ap_done" *)input SEIDEL2D_4__ap_done;
  (* RS_FF = "SEIDEL2D_4__ap_idle" *)input SEIDEL2D_4__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_5.ap_start" *)output SEIDEL2D_5__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_5.ap_ready" *)input SEIDEL2D_5__ap_ready;
  (* RS_FF = "SEIDEL2D_5__ap_done" *)input SEIDEL2D_5__ap_done;
  (* RS_FF = "SEIDEL2D_5__ap_idle" *)input SEIDEL2D_5__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_6.ap_start" *)output SEIDEL2D_6__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_6.ap_ready" *)input SEIDEL2D_6__ap_ready;
  (* RS_FF = "SEIDEL2D_6__ap_done" *)input SEIDEL2D_6__ap_done;
  (* RS_FF = "SEIDEL2D_6__ap_idle" *)input SEIDEL2D_6__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_7.ap_start" *)output SEIDEL2D_7__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_7.ap_ready" *)input SEIDEL2D_7__ap_ready;
  (* RS_FF = "SEIDEL2D_7__ap_done" *)input SEIDEL2D_7__ap_done;
  (* RS_FF = "SEIDEL2D_7__ap_idle" *)input SEIDEL2D_7__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_8.ap_start" *)output SEIDEL2D_8__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_8.ap_ready" *)input SEIDEL2D_8__ap_ready;
  (* RS_FF = "SEIDEL2D_8__ap_done" *)input SEIDEL2D_8__ap_done;
  (* RS_FF = "SEIDEL2D_8__ap_idle" *)input SEIDEL2D_8__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_9.ap_start" *)output SEIDEL2D_9__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_9.ap_ready" *)input SEIDEL2D_9__ap_ready;
  (* RS_FF = "SEIDEL2D_9__ap_done" *)input SEIDEL2D_9__ap_done;
  (* RS_FF = "SEIDEL2D_9__ap_idle" *)input SEIDEL2D_9__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_10.ap_start" *)output SEIDEL2D_10__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_10.ap_ready" *)input SEIDEL2D_10__ap_ready;
  (* RS_FF = "SEIDEL2D_10__ap_done" *)input SEIDEL2D_10__ap_done;
  (* RS_FF = "SEIDEL2D_10__ap_idle" *)input SEIDEL2D_10__ap_idle;
  (* RS_AP_CTRL = "SEIDEL2D_11.ap_start" *)output SEIDEL2D_11__ap_start;
  (* RS_AP_CTRL = "SEIDEL2D_11.ap_ready" *)input SEIDEL2D_11__ap_ready;
  (* RS_FF = "SEIDEL2D_11__ap_done" *)input SEIDEL2D_11__ap_done;
  (* RS_FF = "SEIDEL2D_11__ap_idle" *)input SEIDEL2D_11__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_0.ap_start" *)output inter_kernel_0__ap_start;
  (* RS_AP_CTRL = "inter_kernel_0.ap_ready" *)input inter_kernel_0__ap_ready;
  (* RS_FF = "inter_kernel_0__ap_done" *)input inter_kernel_0__ap_done;
  (* RS_FF = "inter_kernel_0__ap_idle" *)input inter_kernel_0__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_1.ap_start" *)output inter_kernel_1__ap_start;
  (* RS_AP_CTRL = "inter_kernel_1.ap_ready" *)input inter_kernel_1__ap_ready;
  (* RS_FF = "inter_kernel_1__ap_done" *)input inter_kernel_1__ap_done;
  (* RS_FF = "inter_kernel_1__ap_idle" *)input inter_kernel_1__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_2.ap_start" *)output inter_kernel_2__ap_start;
  (* RS_AP_CTRL = "inter_kernel_2.ap_ready" *)input inter_kernel_2__ap_ready;
  (* RS_FF = "inter_kernel_2__ap_done" *)input inter_kernel_2__ap_done;
  (* RS_FF = "inter_kernel_2__ap_idle" *)input inter_kernel_2__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_3.ap_start" *)output inter_kernel_3__ap_start;
  (* RS_AP_CTRL = "inter_kernel_3.ap_ready" *)input inter_kernel_3__ap_ready;
  (* RS_FF = "inter_kernel_3__ap_done" *)input inter_kernel_3__ap_done;
  (* RS_FF = "inter_kernel_3__ap_idle" *)input inter_kernel_3__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_4.ap_start" *)output inter_kernel_4__ap_start;
  (* RS_AP_CTRL = "inter_kernel_4.ap_ready" *)input inter_kernel_4__ap_ready;
  (* RS_FF = "inter_kernel_4__ap_done" *)input inter_kernel_4__ap_done;
  (* RS_FF = "inter_kernel_4__ap_idle" *)input inter_kernel_4__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_5.ap_start" *)output inter_kernel_5__ap_start;
  (* RS_AP_CTRL = "inter_kernel_5.ap_ready" *)input inter_kernel_5__ap_ready;
  (* RS_FF = "inter_kernel_5__ap_done" *)input inter_kernel_5__ap_done;
  (* RS_FF = "inter_kernel_5__ap_idle" *)input inter_kernel_5__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_6.ap_start" *)output inter_kernel_6__ap_start;
  (* RS_AP_CTRL = "inter_kernel_6.ap_ready" *)input inter_kernel_6__ap_ready;
  (* RS_FF = "inter_kernel_6__ap_done" *)input inter_kernel_6__ap_done;
  (* RS_FF = "inter_kernel_6__ap_idle" *)input inter_kernel_6__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_7.ap_start" *)output inter_kernel_7__ap_start;
  (* RS_AP_CTRL = "inter_kernel_7.ap_ready" *)input inter_kernel_7__ap_ready;
  (* RS_FF = "inter_kernel_7__ap_done" *)input inter_kernel_7__ap_done;
  (* RS_FF = "inter_kernel_7__ap_idle" *)input inter_kernel_7__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_8.ap_start" *)output inter_kernel_8__ap_start;
  (* RS_AP_CTRL = "inter_kernel_8.ap_ready" *)input inter_kernel_8__ap_ready;
  (* RS_FF = "inter_kernel_8__ap_done" *)input inter_kernel_8__ap_done;
  (* RS_FF = "inter_kernel_8__ap_idle" *)input inter_kernel_8__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_9.ap_start" *)output inter_kernel_9__ap_start;
  (* RS_AP_CTRL = "inter_kernel_9.ap_ready" *)input inter_kernel_9__ap_ready;
  (* RS_FF = "inter_kernel_9__ap_done" *)input inter_kernel_9__ap_done;
  (* RS_FF = "inter_kernel_9__ap_idle" *)input inter_kernel_9__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_10.ap_start" *)output inter_kernel_10__ap_start;
  (* RS_AP_CTRL = "inter_kernel_10.ap_ready" *)input inter_kernel_10__ap_ready;
  (* RS_FF = "inter_kernel_10__ap_done" *)input inter_kernel_10__ap_done;
  (* RS_FF = "inter_kernel_10__ap_idle" *)input inter_kernel_10__ap_idle;
  (* RS_AP_CTRL = "inter_kernel_11.ap_start" *)output inter_kernel_11__ap_start;
  (* RS_AP_CTRL = "inter_kernel_11.ap_ready" *)input inter_kernel_11__ap_ready;
  (* RS_FF = "inter_kernel_11__ap_done" *)input inter_kernel_11__ap_done;
  (* RS_FF = "inter_kernel_11__ap_idle" *)input inter_kernel_11__ap_idle;
  wire SEIDEL2D_0__ap_start_global__q0;
  wire SEIDEL2D_0__is_done__q0;
  wire SEIDEL2D_0__ap_done_global__q0;
  wire SEIDEL2D_0__ap_start;
  wire SEIDEL2D_0__ap_ready;
  wire SEIDEL2D_0__ap_done;
  wire SEIDEL2D_0__ap_idle;
  reg [1:0] SEIDEL2D_0__state;
  wire SEIDEL2D_1__ap_start_global__q0;
  wire SEIDEL2D_1__is_done__q0;
  wire SEIDEL2D_1__ap_done_global__q0;
  wire SEIDEL2D_1__ap_start;
  wire SEIDEL2D_1__ap_ready;
  wire SEIDEL2D_1__ap_done;
  wire SEIDEL2D_1__ap_idle;
  reg [1:0] SEIDEL2D_1__state;
  wire SEIDEL2D_2__ap_start_global__q0;
  wire SEIDEL2D_2__is_done__q0;
  wire SEIDEL2D_2__ap_done_global__q0;
  wire SEIDEL2D_2__ap_start;
  wire SEIDEL2D_2__ap_ready;
  wire SEIDEL2D_2__ap_done;
  wire SEIDEL2D_2__ap_idle;
  reg [1:0] SEIDEL2D_2__state;
  wire SEIDEL2D_3__ap_start_global__q0;
  wire SEIDEL2D_3__is_done__q0;
  wire SEIDEL2D_3__ap_done_global__q0;
  wire SEIDEL2D_3__ap_start;
  wire SEIDEL2D_3__ap_ready;
  wire SEIDEL2D_3__ap_done;
  wire SEIDEL2D_3__ap_idle;
  reg [1:0] SEIDEL2D_3__state;
  wire SEIDEL2D_4__ap_start_global__q0;
  wire SEIDEL2D_4__is_done__q0;
  wire SEIDEL2D_4__ap_done_global__q0;
  wire SEIDEL2D_4__ap_start;
  wire SEIDEL2D_4__ap_ready;
  wire SEIDEL2D_4__ap_done;
  wire SEIDEL2D_4__ap_idle;
  reg [1:0] SEIDEL2D_4__state;
  wire SEIDEL2D_5__ap_start_global__q0;
  wire SEIDEL2D_5__is_done__q0;
  wire SEIDEL2D_5__ap_done_global__q0;
  wire SEIDEL2D_5__ap_start;
  wire SEIDEL2D_5__ap_ready;
  wire SEIDEL2D_5__ap_done;
  wire SEIDEL2D_5__ap_idle;
  reg [1:0] SEIDEL2D_5__state;
  wire SEIDEL2D_6__ap_start_global__q0;
  wire SEIDEL2D_6__is_done__q0;
  wire SEIDEL2D_6__ap_done_global__q0;
  wire SEIDEL2D_6__ap_start;
  wire SEIDEL2D_6__ap_ready;
  wire SEIDEL2D_6__ap_done;
  wire SEIDEL2D_6__ap_idle;
  reg [1:0] SEIDEL2D_6__state;
  wire SEIDEL2D_7__ap_start_global__q0;
  wire SEIDEL2D_7__is_done__q0;
  wire SEIDEL2D_7__ap_done_global__q0;
  wire SEIDEL2D_7__ap_start;
  wire SEIDEL2D_7__ap_ready;
  wire SEIDEL2D_7__ap_done;
  wire SEIDEL2D_7__ap_idle;
  reg [1:0] SEIDEL2D_7__state;
  wire SEIDEL2D_8__ap_start_global__q0;
  wire SEIDEL2D_8__is_done__q0;
  wire SEIDEL2D_8__ap_done_global__q0;
  wire SEIDEL2D_8__ap_start;
  wire SEIDEL2D_8__ap_ready;
  wire SEIDEL2D_8__ap_done;
  wire SEIDEL2D_8__ap_idle;
  reg [1:0] SEIDEL2D_8__state;
  wire SEIDEL2D_9__ap_start_global__q0;
  wire SEIDEL2D_9__is_done__q0;
  wire SEIDEL2D_9__ap_done_global__q0;
  wire SEIDEL2D_9__ap_start;
  wire SEIDEL2D_9__ap_ready;
  wire SEIDEL2D_9__ap_done;
  wire SEIDEL2D_9__ap_idle;
  reg [1:0] SEIDEL2D_9__state;
  wire SEIDEL2D_10__ap_start_global__q0;
  wire SEIDEL2D_10__is_done__q0;
  wire SEIDEL2D_10__ap_done_global__q0;
  wire SEIDEL2D_10__ap_start;
  wire SEIDEL2D_10__ap_ready;
  wire SEIDEL2D_10__ap_done;
  wire SEIDEL2D_10__ap_idle;
  reg [1:0] SEIDEL2D_10__state;
  wire SEIDEL2D_11__ap_start_global__q0;
  wire SEIDEL2D_11__is_done__q0;
  wire SEIDEL2D_11__ap_done_global__q0;
  wire SEIDEL2D_11__ap_start;
  wire SEIDEL2D_11__ap_ready;
  wire SEIDEL2D_11__ap_done;
  wire SEIDEL2D_11__ap_idle;
  reg [1:0] SEIDEL2D_11__state;
  wire inter_kernel_0__ap_start_global__q0;
  wire inter_kernel_0__is_done__q0;
  wire inter_kernel_0__ap_done_global__q0;
  wire inter_kernel_0__ap_start;
  wire inter_kernel_0__ap_ready;
  wire inter_kernel_0__ap_done;
  wire inter_kernel_0__ap_idle;
  reg [1:0] inter_kernel_0__state;
  wire inter_kernel_1__ap_start_global__q0;
  wire inter_kernel_1__is_done__q0;
  wire inter_kernel_1__ap_done_global__q0;
  wire inter_kernel_1__ap_start;
  wire inter_kernel_1__ap_ready;
  wire inter_kernel_1__ap_done;
  wire inter_kernel_1__ap_idle;
  reg [1:0] inter_kernel_1__state;
  wire inter_kernel_2__ap_start_global__q0;
  wire inter_kernel_2__is_done__q0;
  wire inter_kernel_2__ap_done_global__q0;
  wire inter_kernel_2__ap_start;
  wire inter_kernel_2__ap_ready;
  wire inter_kernel_2__ap_done;
  wire inter_kernel_2__ap_idle;
  reg [1:0] inter_kernel_2__state;
  wire inter_kernel_3__ap_start_global__q0;
  wire inter_kernel_3__is_done__q0;
  wire inter_kernel_3__ap_done_global__q0;
  wire inter_kernel_3__ap_start;
  wire inter_kernel_3__ap_ready;
  wire inter_kernel_3__ap_done;
  wire inter_kernel_3__ap_idle;
  reg [1:0] inter_kernel_3__state;
  wire inter_kernel_4__ap_start_global__q0;
  wire inter_kernel_4__is_done__q0;
  wire inter_kernel_4__ap_done_global__q0;
  wire inter_kernel_4__ap_start;
  wire inter_kernel_4__ap_ready;
  wire inter_kernel_4__ap_done;
  wire inter_kernel_4__ap_idle;
  reg [1:0] inter_kernel_4__state;
  wire inter_kernel_5__ap_start_global__q0;
  wire inter_kernel_5__is_done__q0;
  wire inter_kernel_5__ap_done_global__q0;
  wire inter_kernel_5__ap_start;
  wire inter_kernel_5__ap_ready;
  wire inter_kernel_5__ap_done;
  wire inter_kernel_5__ap_idle;
  reg [1:0] inter_kernel_5__state;
  wire inter_kernel_6__ap_start_global__q0;
  wire inter_kernel_6__is_done__q0;
  wire inter_kernel_6__ap_done_global__q0;
  wire inter_kernel_6__ap_start;
  wire inter_kernel_6__ap_ready;
  wire inter_kernel_6__ap_done;
  wire inter_kernel_6__ap_idle;
  reg [1:0] inter_kernel_6__state;
  wire inter_kernel_7__ap_start_global__q0;
  wire inter_kernel_7__is_done__q0;
  wire inter_kernel_7__ap_done_global__q0;
  wire inter_kernel_7__ap_start;
  wire inter_kernel_7__ap_ready;
  wire inter_kernel_7__ap_done;
  wire inter_kernel_7__ap_idle;
  reg [1:0] inter_kernel_7__state;
  wire inter_kernel_8__ap_start_global__q0;
  wire inter_kernel_8__is_done__q0;
  wire inter_kernel_8__ap_done_global__q0;
  wire inter_kernel_8__ap_start;
  wire inter_kernel_8__ap_ready;
  wire inter_kernel_8__ap_done;
  wire inter_kernel_8__ap_idle;
  reg [1:0] inter_kernel_8__state;
  wire inter_kernel_9__ap_start_global__q0;
  wire inter_kernel_9__is_done__q0;
  wire inter_kernel_9__ap_done_global__q0;
  wire inter_kernel_9__ap_start;
  wire inter_kernel_9__ap_ready;
  wire inter_kernel_9__ap_done;
  wire inter_kernel_9__ap_idle;
  reg [1:0] inter_kernel_9__state;
  wire inter_kernel_10__ap_start_global__q0;
  wire inter_kernel_10__is_done__q0;
  wire inter_kernel_10__ap_done_global__q0;
  wire inter_kernel_10__ap_start;
  wire inter_kernel_10__ap_ready;
  wire inter_kernel_10__ap_done;
  wire inter_kernel_10__ap_idle;
  reg [1:0] inter_kernel_10__state;
  wire inter_kernel_11__ap_start_global__q0;
  wire inter_kernel_11__is_done__q0;
  wire inter_kernel_11__ap_done_global__q0;
  wire inter_kernel_11__ap_start;
  wire inter_kernel_11__ap_ready;
  wire inter_kernel_11__ap_done;
  wire inter_kernel_11__ap_idle;
  reg [1:0] inter_kernel_11__state;
  reg [1:0] tapa_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  wire ap_done__q0;
  assign SEIDEL2D_0__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_0__is_done__q0 = (SEIDEL2D_0__state == 2'b10);
  assign SEIDEL2D_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_0__state <= 2'b00;
    end else begin
      if(SEIDEL2D_0__state == 2'b00) begin
        if(SEIDEL2D_0__ap_start_global__q0) begin
          SEIDEL2D_0__state <= 2'b01;
        end
      end
      if(SEIDEL2D_0__state == 2'b01) begin
        if(SEIDEL2D_0__ap_ready) begin
          if(SEIDEL2D_0__ap_done) begin
            SEIDEL2D_0__state <= 2'b10;
          end else begin
            SEIDEL2D_0__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_0__state == 2'b11) begin
        if(SEIDEL2D_0__ap_done) begin
          SEIDEL2D_0__state <= 2'b10;
        end
      end
      if(SEIDEL2D_0__state == 2'b10) begin
        if(SEIDEL2D_0__ap_done_global__q0) begin
          SEIDEL2D_0__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_0__ap_start = (SEIDEL2D_0__state == 2'b01);
  assign SEIDEL2D_1__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_1__is_done__q0 = (SEIDEL2D_1__state == 2'b10);
  assign SEIDEL2D_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_1__state <= 2'b00;
    end else begin
      if(SEIDEL2D_1__state == 2'b00) begin
        if(SEIDEL2D_1__ap_start_global__q0) begin
          SEIDEL2D_1__state <= 2'b01;
        end
      end
      if(SEIDEL2D_1__state == 2'b01) begin
        if(SEIDEL2D_1__ap_ready) begin
          if(SEIDEL2D_1__ap_done) begin
            SEIDEL2D_1__state <= 2'b10;
          end else begin
            SEIDEL2D_1__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_1__state == 2'b11) begin
        if(SEIDEL2D_1__ap_done) begin
          SEIDEL2D_1__state <= 2'b10;
        end
      end
      if(SEIDEL2D_1__state == 2'b10) begin
        if(SEIDEL2D_1__ap_done_global__q0) begin
          SEIDEL2D_1__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_1__ap_start = (SEIDEL2D_1__state == 2'b01);
  assign SEIDEL2D_2__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_2__is_done__q0 = (SEIDEL2D_2__state == 2'b10);
  assign SEIDEL2D_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_2__state <= 2'b00;
    end else begin
      if(SEIDEL2D_2__state == 2'b00) begin
        if(SEIDEL2D_2__ap_start_global__q0) begin
          SEIDEL2D_2__state <= 2'b01;
        end
      end
      if(SEIDEL2D_2__state == 2'b01) begin
        if(SEIDEL2D_2__ap_ready) begin
          if(SEIDEL2D_2__ap_done) begin
            SEIDEL2D_2__state <= 2'b10;
          end else begin
            SEIDEL2D_2__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_2__state == 2'b11) begin
        if(SEIDEL2D_2__ap_done) begin
          SEIDEL2D_2__state <= 2'b10;
        end
      end
      if(SEIDEL2D_2__state == 2'b10) begin
        if(SEIDEL2D_2__ap_done_global__q0) begin
          SEIDEL2D_2__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_2__ap_start = (SEIDEL2D_2__state == 2'b01);
  assign SEIDEL2D_3__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_3__is_done__q0 = (SEIDEL2D_3__state == 2'b10);
  assign SEIDEL2D_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_3__state <= 2'b00;
    end else begin
      if(SEIDEL2D_3__state == 2'b00) begin
        if(SEIDEL2D_3__ap_start_global__q0) begin
          SEIDEL2D_3__state <= 2'b01;
        end
      end
      if(SEIDEL2D_3__state == 2'b01) begin
        if(SEIDEL2D_3__ap_ready) begin
          if(SEIDEL2D_3__ap_done) begin
            SEIDEL2D_3__state <= 2'b10;
          end else begin
            SEIDEL2D_3__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_3__state == 2'b11) begin
        if(SEIDEL2D_3__ap_done) begin
          SEIDEL2D_3__state <= 2'b10;
        end
      end
      if(SEIDEL2D_3__state == 2'b10) begin
        if(SEIDEL2D_3__ap_done_global__q0) begin
          SEIDEL2D_3__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_3__ap_start = (SEIDEL2D_3__state == 2'b01);
  assign SEIDEL2D_4__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_4__is_done__q0 = (SEIDEL2D_4__state == 2'b10);
  assign SEIDEL2D_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_4__state <= 2'b00;
    end else begin
      if(SEIDEL2D_4__state == 2'b00) begin
        if(SEIDEL2D_4__ap_start_global__q0) begin
          SEIDEL2D_4__state <= 2'b01;
        end
      end
      if(SEIDEL2D_4__state == 2'b01) begin
        if(SEIDEL2D_4__ap_ready) begin
          if(SEIDEL2D_4__ap_done) begin
            SEIDEL2D_4__state <= 2'b10;
          end else begin
            SEIDEL2D_4__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_4__state == 2'b11) begin
        if(SEIDEL2D_4__ap_done) begin
          SEIDEL2D_4__state <= 2'b10;
        end
      end
      if(SEIDEL2D_4__state == 2'b10) begin
        if(SEIDEL2D_4__ap_done_global__q0) begin
          SEIDEL2D_4__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_4__ap_start = (SEIDEL2D_4__state == 2'b01);
  assign SEIDEL2D_5__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_5__is_done__q0 = (SEIDEL2D_5__state == 2'b10);
  assign SEIDEL2D_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_5__state <= 2'b00;
    end else begin
      if(SEIDEL2D_5__state == 2'b00) begin
        if(SEIDEL2D_5__ap_start_global__q0) begin
          SEIDEL2D_5__state <= 2'b01;
        end
      end
      if(SEIDEL2D_5__state == 2'b01) begin
        if(SEIDEL2D_5__ap_ready) begin
          if(SEIDEL2D_5__ap_done) begin
            SEIDEL2D_5__state <= 2'b10;
          end else begin
            SEIDEL2D_5__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_5__state == 2'b11) begin
        if(SEIDEL2D_5__ap_done) begin
          SEIDEL2D_5__state <= 2'b10;
        end
      end
      if(SEIDEL2D_5__state == 2'b10) begin
        if(SEIDEL2D_5__ap_done_global__q0) begin
          SEIDEL2D_5__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_5__ap_start = (SEIDEL2D_5__state == 2'b01);
  assign SEIDEL2D_6__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_6__is_done__q0 = (SEIDEL2D_6__state == 2'b10);
  assign SEIDEL2D_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_6__state <= 2'b00;
    end else begin
      if(SEIDEL2D_6__state == 2'b00) begin
        if(SEIDEL2D_6__ap_start_global__q0) begin
          SEIDEL2D_6__state <= 2'b01;
        end
      end
      if(SEIDEL2D_6__state == 2'b01) begin
        if(SEIDEL2D_6__ap_ready) begin
          if(SEIDEL2D_6__ap_done) begin
            SEIDEL2D_6__state <= 2'b10;
          end else begin
            SEIDEL2D_6__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_6__state == 2'b11) begin
        if(SEIDEL2D_6__ap_done) begin
          SEIDEL2D_6__state <= 2'b10;
        end
      end
      if(SEIDEL2D_6__state == 2'b10) begin
        if(SEIDEL2D_6__ap_done_global__q0) begin
          SEIDEL2D_6__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_6__ap_start = (SEIDEL2D_6__state == 2'b01);
  assign SEIDEL2D_7__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_7__is_done__q0 = (SEIDEL2D_7__state == 2'b10);
  assign SEIDEL2D_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_7__state <= 2'b00;
    end else begin
      if(SEIDEL2D_7__state == 2'b00) begin
        if(SEIDEL2D_7__ap_start_global__q0) begin
          SEIDEL2D_7__state <= 2'b01;
        end
      end
      if(SEIDEL2D_7__state == 2'b01) begin
        if(SEIDEL2D_7__ap_ready) begin
          if(SEIDEL2D_7__ap_done) begin
            SEIDEL2D_7__state <= 2'b10;
          end else begin
            SEIDEL2D_7__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_7__state == 2'b11) begin
        if(SEIDEL2D_7__ap_done) begin
          SEIDEL2D_7__state <= 2'b10;
        end
      end
      if(SEIDEL2D_7__state == 2'b10) begin
        if(SEIDEL2D_7__ap_done_global__q0) begin
          SEIDEL2D_7__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_7__ap_start = (SEIDEL2D_7__state == 2'b01);
  assign SEIDEL2D_8__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_8__is_done__q0 = (SEIDEL2D_8__state == 2'b10);
  assign SEIDEL2D_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_8__state <= 2'b00;
    end else begin
      if(SEIDEL2D_8__state == 2'b00) begin
        if(SEIDEL2D_8__ap_start_global__q0) begin
          SEIDEL2D_8__state <= 2'b01;
        end
      end
      if(SEIDEL2D_8__state == 2'b01) begin
        if(SEIDEL2D_8__ap_ready) begin
          if(SEIDEL2D_8__ap_done) begin
            SEIDEL2D_8__state <= 2'b10;
          end else begin
            SEIDEL2D_8__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_8__state == 2'b11) begin
        if(SEIDEL2D_8__ap_done) begin
          SEIDEL2D_8__state <= 2'b10;
        end
      end
      if(SEIDEL2D_8__state == 2'b10) begin
        if(SEIDEL2D_8__ap_done_global__q0) begin
          SEIDEL2D_8__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_8__ap_start = (SEIDEL2D_8__state == 2'b01);
  assign SEIDEL2D_9__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_9__is_done__q0 = (SEIDEL2D_9__state == 2'b10);
  assign SEIDEL2D_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_9__state <= 2'b00;
    end else begin
      if(SEIDEL2D_9__state == 2'b00) begin
        if(SEIDEL2D_9__ap_start_global__q0) begin
          SEIDEL2D_9__state <= 2'b01;
        end
      end
      if(SEIDEL2D_9__state == 2'b01) begin
        if(SEIDEL2D_9__ap_ready) begin
          if(SEIDEL2D_9__ap_done) begin
            SEIDEL2D_9__state <= 2'b10;
          end else begin
            SEIDEL2D_9__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_9__state == 2'b11) begin
        if(SEIDEL2D_9__ap_done) begin
          SEIDEL2D_9__state <= 2'b10;
        end
      end
      if(SEIDEL2D_9__state == 2'b10) begin
        if(SEIDEL2D_9__ap_done_global__q0) begin
          SEIDEL2D_9__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_9__ap_start = (SEIDEL2D_9__state == 2'b01);
  assign SEIDEL2D_10__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_10__is_done__q0 = (SEIDEL2D_10__state == 2'b10);
  assign SEIDEL2D_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_10__state <= 2'b00;
    end else begin
      if(SEIDEL2D_10__state == 2'b00) begin
        if(SEIDEL2D_10__ap_start_global__q0) begin
          SEIDEL2D_10__state <= 2'b01;
        end
      end
      if(SEIDEL2D_10__state == 2'b01) begin
        if(SEIDEL2D_10__ap_ready) begin
          if(SEIDEL2D_10__ap_done) begin
            SEIDEL2D_10__state <= 2'b10;
          end else begin
            SEIDEL2D_10__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_10__state == 2'b11) begin
        if(SEIDEL2D_10__ap_done) begin
          SEIDEL2D_10__state <= 2'b10;
        end
      end
      if(SEIDEL2D_10__state == 2'b10) begin
        if(SEIDEL2D_10__ap_done_global__q0) begin
          SEIDEL2D_10__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_10__ap_start = (SEIDEL2D_10__state == 2'b01);
  assign SEIDEL2D_11__ap_start_global__q0 = ap_start__q0;
  assign SEIDEL2D_11__is_done__q0 = (SEIDEL2D_11__state == 2'b10);
  assign SEIDEL2D_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      SEIDEL2D_11__state <= 2'b00;
    end else begin
      if(SEIDEL2D_11__state == 2'b00) begin
        if(SEIDEL2D_11__ap_start_global__q0) begin
          SEIDEL2D_11__state <= 2'b01;
        end
      end
      if(SEIDEL2D_11__state == 2'b01) begin
        if(SEIDEL2D_11__ap_ready) begin
          if(SEIDEL2D_11__ap_done) begin
            SEIDEL2D_11__state <= 2'b10;
          end else begin
            SEIDEL2D_11__state <= 2'b11;
          end
        end
      end
      if(SEIDEL2D_11__state == 2'b11) begin
        if(SEIDEL2D_11__ap_done) begin
          SEIDEL2D_11__state <= 2'b10;
        end
      end
      if(SEIDEL2D_11__state == 2'b10) begin
        if(SEIDEL2D_11__ap_done_global__q0) begin
          SEIDEL2D_11__state <= 2'b00;
        end
      end
    end
  end

  assign SEIDEL2D_11__ap_start = (SEIDEL2D_11__state == 2'b01);
  assign inter_kernel_0__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_0__is_done__q0 = (inter_kernel_0__state == 2'b10);
  assign inter_kernel_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_0__state <= 2'b00;
    end else begin
      if(inter_kernel_0__state == 2'b00) begin
        if(inter_kernel_0__ap_start_global__q0) begin
          inter_kernel_0__state <= 2'b01;
        end
      end
      if(inter_kernel_0__state == 2'b01) begin
        if(inter_kernel_0__ap_ready) begin
          if(inter_kernel_0__ap_done) begin
            inter_kernel_0__state <= 2'b10;
          end else begin
            inter_kernel_0__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_0__state == 2'b11) begin
        if(inter_kernel_0__ap_done) begin
          inter_kernel_0__state <= 2'b10;
        end
      end
      if(inter_kernel_0__state == 2'b10) begin
        if(inter_kernel_0__ap_done_global__q0) begin
          inter_kernel_0__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_0__ap_start = (inter_kernel_0__state == 2'b01);
  assign inter_kernel_1__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_1__is_done__q0 = (inter_kernel_1__state == 2'b10);
  assign inter_kernel_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_1__state <= 2'b00;
    end else begin
      if(inter_kernel_1__state == 2'b00) begin
        if(inter_kernel_1__ap_start_global__q0) begin
          inter_kernel_1__state <= 2'b01;
        end
      end
      if(inter_kernel_1__state == 2'b01) begin
        if(inter_kernel_1__ap_ready) begin
          if(inter_kernel_1__ap_done) begin
            inter_kernel_1__state <= 2'b10;
          end else begin
            inter_kernel_1__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_1__state == 2'b11) begin
        if(inter_kernel_1__ap_done) begin
          inter_kernel_1__state <= 2'b10;
        end
      end
      if(inter_kernel_1__state == 2'b10) begin
        if(inter_kernel_1__ap_done_global__q0) begin
          inter_kernel_1__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_1__ap_start = (inter_kernel_1__state == 2'b01);
  assign inter_kernel_2__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_2__is_done__q0 = (inter_kernel_2__state == 2'b10);
  assign inter_kernel_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_2__state <= 2'b00;
    end else begin
      if(inter_kernel_2__state == 2'b00) begin
        if(inter_kernel_2__ap_start_global__q0) begin
          inter_kernel_2__state <= 2'b01;
        end
      end
      if(inter_kernel_2__state == 2'b01) begin
        if(inter_kernel_2__ap_ready) begin
          if(inter_kernel_2__ap_done) begin
            inter_kernel_2__state <= 2'b10;
          end else begin
            inter_kernel_2__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_2__state == 2'b11) begin
        if(inter_kernel_2__ap_done) begin
          inter_kernel_2__state <= 2'b10;
        end
      end
      if(inter_kernel_2__state == 2'b10) begin
        if(inter_kernel_2__ap_done_global__q0) begin
          inter_kernel_2__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_2__ap_start = (inter_kernel_2__state == 2'b01);
  assign inter_kernel_3__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_3__is_done__q0 = (inter_kernel_3__state == 2'b10);
  assign inter_kernel_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_3__state <= 2'b00;
    end else begin
      if(inter_kernel_3__state == 2'b00) begin
        if(inter_kernel_3__ap_start_global__q0) begin
          inter_kernel_3__state <= 2'b01;
        end
      end
      if(inter_kernel_3__state == 2'b01) begin
        if(inter_kernel_3__ap_ready) begin
          if(inter_kernel_3__ap_done) begin
            inter_kernel_3__state <= 2'b10;
          end else begin
            inter_kernel_3__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_3__state == 2'b11) begin
        if(inter_kernel_3__ap_done) begin
          inter_kernel_3__state <= 2'b10;
        end
      end
      if(inter_kernel_3__state == 2'b10) begin
        if(inter_kernel_3__ap_done_global__q0) begin
          inter_kernel_3__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_3__ap_start = (inter_kernel_3__state == 2'b01);
  assign inter_kernel_4__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_4__is_done__q0 = (inter_kernel_4__state == 2'b10);
  assign inter_kernel_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_4__state <= 2'b00;
    end else begin
      if(inter_kernel_4__state == 2'b00) begin
        if(inter_kernel_4__ap_start_global__q0) begin
          inter_kernel_4__state <= 2'b01;
        end
      end
      if(inter_kernel_4__state == 2'b01) begin
        if(inter_kernel_4__ap_ready) begin
          if(inter_kernel_4__ap_done) begin
            inter_kernel_4__state <= 2'b10;
          end else begin
            inter_kernel_4__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_4__state == 2'b11) begin
        if(inter_kernel_4__ap_done) begin
          inter_kernel_4__state <= 2'b10;
        end
      end
      if(inter_kernel_4__state == 2'b10) begin
        if(inter_kernel_4__ap_done_global__q0) begin
          inter_kernel_4__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_4__ap_start = (inter_kernel_4__state == 2'b01);
  assign inter_kernel_5__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_5__is_done__q0 = (inter_kernel_5__state == 2'b10);
  assign inter_kernel_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_5__state <= 2'b00;
    end else begin
      if(inter_kernel_5__state == 2'b00) begin
        if(inter_kernel_5__ap_start_global__q0) begin
          inter_kernel_5__state <= 2'b01;
        end
      end
      if(inter_kernel_5__state == 2'b01) begin
        if(inter_kernel_5__ap_ready) begin
          if(inter_kernel_5__ap_done) begin
            inter_kernel_5__state <= 2'b10;
          end else begin
            inter_kernel_5__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_5__state == 2'b11) begin
        if(inter_kernel_5__ap_done) begin
          inter_kernel_5__state <= 2'b10;
        end
      end
      if(inter_kernel_5__state == 2'b10) begin
        if(inter_kernel_5__ap_done_global__q0) begin
          inter_kernel_5__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_5__ap_start = (inter_kernel_5__state == 2'b01);
  assign inter_kernel_6__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_6__is_done__q0 = (inter_kernel_6__state == 2'b10);
  assign inter_kernel_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_6__state <= 2'b00;
    end else begin
      if(inter_kernel_6__state == 2'b00) begin
        if(inter_kernel_6__ap_start_global__q0) begin
          inter_kernel_6__state <= 2'b01;
        end
      end
      if(inter_kernel_6__state == 2'b01) begin
        if(inter_kernel_6__ap_ready) begin
          if(inter_kernel_6__ap_done) begin
            inter_kernel_6__state <= 2'b10;
          end else begin
            inter_kernel_6__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_6__state == 2'b11) begin
        if(inter_kernel_6__ap_done) begin
          inter_kernel_6__state <= 2'b10;
        end
      end
      if(inter_kernel_6__state == 2'b10) begin
        if(inter_kernel_6__ap_done_global__q0) begin
          inter_kernel_6__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_6__ap_start = (inter_kernel_6__state == 2'b01);
  assign inter_kernel_7__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_7__is_done__q0 = (inter_kernel_7__state == 2'b10);
  assign inter_kernel_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_7__state <= 2'b00;
    end else begin
      if(inter_kernel_7__state == 2'b00) begin
        if(inter_kernel_7__ap_start_global__q0) begin
          inter_kernel_7__state <= 2'b01;
        end
      end
      if(inter_kernel_7__state == 2'b01) begin
        if(inter_kernel_7__ap_ready) begin
          if(inter_kernel_7__ap_done) begin
            inter_kernel_7__state <= 2'b10;
          end else begin
            inter_kernel_7__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_7__state == 2'b11) begin
        if(inter_kernel_7__ap_done) begin
          inter_kernel_7__state <= 2'b10;
        end
      end
      if(inter_kernel_7__state == 2'b10) begin
        if(inter_kernel_7__ap_done_global__q0) begin
          inter_kernel_7__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_7__ap_start = (inter_kernel_7__state == 2'b01);
  assign inter_kernel_8__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_8__is_done__q0 = (inter_kernel_8__state == 2'b10);
  assign inter_kernel_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_8__state <= 2'b00;
    end else begin
      if(inter_kernel_8__state == 2'b00) begin
        if(inter_kernel_8__ap_start_global__q0) begin
          inter_kernel_8__state <= 2'b01;
        end
      end
      if(inter_kernel_8__state == 2'b01) begin
        if(inter_kernel_8__ap_ready) begin
          if(inter_kernel_8__ap_done) begin
            inter_kernel_8__state <= 2'b10;
          end else begin
            inter_kernel_8__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_8__state == 2'b11) begin
        if(inter_kernel_8__ap_done) begin
          inter_kernel_8__state <= 2'b10;
        end
      end
      if(inter_kernel_8__state == 2'b10) begin
        if(inter_kernel_8__ap_done_global__q0) begin
          inter_kernel_8__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_8__ap_start = (inter_kernel_8__state == 2'b01);
  assign inter_kernel_9__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_9__is_done__q0 = (inter_kernel_9__state == 2'b10);
  assign inter_kernel_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_9__state <= 2'b00;
    end else begin
      if(inter_kernel_9__state == 2'b00) begin
        if(inter_kernel_9__ap_start_global__q0) begin
          inter_kernel_9__state <= 2'b01;
        end
      end
      if(inter_kernel_9__state == 2'b01) begin
        if(inter_kernel_9__ap_ready) begin
          if(inter_kernel_9__ap_done) begin
            inter_kernel_9__state <= 2'b10;
          end else begin
            inter_kernel_9__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_9__state == 2'b11) begin
        if(inter_kernel_9__ap_done) begin
          inter_kernel_9__state <= 2'b10;
        end
      end
      if(inter_kernel_9__state == 2'b10) begin
        if(inter_kernel_9__ap_done_global__q0) begin
          inter_kernel_9__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_9__ap_start = (inter_kernel_9__state == 2'b01);
  assign inter_kernel_10__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_10__is_done__q0 = (inter_kernel_10__state == 2'b10);
  assign inter_kernel_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_10__state <= 2'b00;
    end else begin
      if(inter_kernel_10__state == 2'b00) begin
        if(inter_kernel_10__ap_start_global__q0) begin
          inter_kernel_10__state <= 2'b01;
        end
      end
      if(inter_kernel_10__state == 2'b01) begin
        if(inter_kernel_10__ap_ready) begin
          if(inter_kernel_10__ap_done) begin
            inter_kernel_10__state <= 2'b10;
          end else begin
            inter_kernel_10__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_10__state == 2'b11) begin
        if(inter_kernel_10__ap_done) begin
          inter_kernel_10__state <= 2'b10;
        end
      end
      if(inter_kernel_10__state == 2'b10) begin
        if(inter_kernel_10__ap_done_global__q0) begin
          inter_kernel_10__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_10__ap_start = (inter_kernel_10__state == 2'b01);
  assign inter_kernel_11__ap_start_global__q0 = ap_start__q0;
  assign inter_kernel_11__is_done__q0 = (inter_kernel_11__state == 2'b10);
  assign inter_kernel_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      inter_kernel_11__state <= 2'b00;
    end else begin
      if(inter_kernel_11__state == 2'b00) begin
        if(inter_kernel_11__ap_start_global__q0) begin
          inter_kernel_11__state <= 2'b01;
        end
      end
      if(inter_kernel_11__state == 2'b01) begin
        if(inter_kernel_11__ap_ready) begin
          if(inter_kernel_11__ap_done) begin
            inter_kernel_11__state <= 2'b10;
          end else begin
            inter_kernel_11__state <= 2'b11;
          end
        end
      end
      if(inter_kernel_11__state == 2'b11) begin
        if(inter_kernel_11__ap_done) begin
          inter_kernel_11__state <= 2'b10;
        end
      end
      if(inter_kernel_11__state == 2'b10) begin
        if(inter_kernel_11__ap_done_global__q0) begin
          inter_kernel_11__state <= 2'b00;
        end
      end
    end
  end

  assign inter_kernel_11__ap_start = (inter_kernel_11__state == 2'b01);

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      tapa_state <= 2'b00;
    end else begin
      case(tapa_state)
        2'b00: begin
          if(ap_start__q0) begin
            tapa_state <= 2'b01;
          end
        end
        2'b01: begin
          if(SEIDEL2D_0__is_done__q0 && SEIDEL2D_1__is_done__q0 && SEIDEL2D_2__is_done__q0 && SEIDEL2D_3__is_done__q0 && SEIDEL2D_4__is_done__q0 && SEIDEL2D_5__is_done__q0 && SEIDEL2D_6__is_done__q0 && SEIDEL2D_7__is_done__q0 && SEIDEL2D_8__is_done__q0 && SEIDEL2D_9__is_done__q0 && SEIDEL2D_10__is_done__q0 && SEIDEL2D_11__is_done__q0 && inter_kernel_0__is_done__q0 && inter_kernel_1__is_done__q0 && inter_kernel_2__is_done__q0 && inter_kernel_3__is_done__q0 && inter_kernel_4__is_done__q0 && inter_kernel_5__is_done__q0 && inter_kernel_6__is_done__q0 && inter_kernel_7__is_done__q0 && inter_kernel_8__is_done__q0 && inter_kernel_9__is_done__q0 && inter_kernel_10__is_done__q0 && inter_kernel_11__is_done__q0) begin
            tapa_state <= 2'b10;
          end
        end
        2'b10: begin
          tapa_state <= 2'b00;
          countdown <= 1'd0;
        end
        2'b11: begin
          if(countdown == 1'd0) begin
            tapa_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end
      endcase
    end
  end

  assign ap_idle = (tapa_state == 2'b00);
  assign ap_done = ap_done__q0;
  assign ap_ready = ap_done__q0;
  assign ap_start__q0 = ap_start;
  assign ap_done__q0 = (tapa_state == 2'b10);

endmodule
