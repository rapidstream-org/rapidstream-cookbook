

module vadd_bw_fsm
(
  ap_clk,
  ap_rst_n,
  ap_start,
  ap_ready,
  ap_done,
  ap_idle,
  n,
  rmem0,
  rmem1,
  rmem2,
  rmem3,
  rmem4,
  rmem5,
  rmem6,
  rmem7,
  rmem8,
  rmem9,
  rmem10,
  rmem11,
  rmem12,
  rmem13,
  rmem14,
  rmem15,
  rmem16,
  rmem17,
  rmem18,
  rmem19,
  rmem20,
  rmem21,
  rmem22,
  rmem23,
  rmem24,
  rmem25,
  rmem26,
  rmem27,
  rmem28,
  rmem29,
  wmem0,
  Mmap2Stream_0___n__q0,
  Mmap2Stream_0___rmem0__q0,
  Mmap2Stream_0__ap_start,
  Mmap2Stream_0__ap_ready,
  Mmap2Stream_0__ap_done,
  Mmap2Stream_0__ap_idle,
  Mmap2Stream_1___n__q0,
  Mmap2Stream_1___rmem1__q0,
  Mmap2Stream_1__ap_start,
  Mmap2Stream_1__ap_ready,
  Mmap2Stream_1__ap_done,
  Mmap2Stream_1__ap_idle,
  Mmap2Stream_2___n__q0,
  Mmap2Stream_2___rmem2__q0,
  Mmap2Stream_2__ap_start,
  Mmap2Stream_2__ap_ready,
  Mmap2Stream_2__ap_done,
  Mmap2Stream_2__ap_idle,
  Mmap2Stream_3___n__q0,
  Mmap2Stream_3___rmem3__q0,
  Mmap2Stream_3__ap_start,
  Mmap2Stream_3__ap_ready,
  Mmap2Stream_3__ap_done,
  Mmap2Stream_3__ap_idle,
  Mmap2Stream_4___n__q0,
  Mmap2Stream_4___rmem4__q0,
  Mmap2Stream_4__ap_start,
  Mmap2Stream_4__ap_ready,
  Mmap2Stream_4__ap_done,
  Mmap2Stream_4__ap_idle,
  Mmap2Stream_5___n__q0,
  Mmap2Stream_5___rmem5__q0,
  Mmap2Stream_5__ap_start,
  Mmap2Stream_5__ap_ready,
  Mmap2Stream_5__ap_done,
  Mmap2Stream_5__ap_idle,
  Mmap2Stream_6___n__q0,
  Mmap2Stream_6___rmem6__q0,
  Mmap2Stream_6__ap_start,
  Mmap2Stream_6__ap_ready,
  Mmap2Stream_6__ap_done,
  Mmap2Stream_6__ap_idle,
  Mmap2Stream_7___n__q0,
  Mmap2Stream_7___rmem7__q0,
  Mmap2Stream_7__ap_start,
  Mmap2Stream_7__ap_ready,
  Mmap2Stream_7__ap_done,
  Mmap2Stream_7__ap_idle,
  Mmap2Stream_8___n__q0,
  Mmap2Stream_8___rmem8__q0,
  Mmap2Stream_8__ap_start,
  Mmap2Stream_8__ap_ready,
  Mmap2Stream_8__ap_done,
  Mmap2Stream_8__ap_idle,
  Mmap2Stream_9___n__q0,
  Mmap2Stream_9___rmem9__q0,
  Mmap2Stream_9__ap_start,
  Mmap2Stream_9__ap_ready,
  Mmap2Stream_9__ap_done,
  Mmap2Stream_9__ap_idle,
  Mmap2Stream_10___n__q0,
  Mmap2Stream_10___rmem10__q0,
  Mmap2Stream_10__ap_start,
  Mmap2Stream_10__ap_ready,
  Mmap2Stream_10__ap_done,
  Mmap2Stream_10__ap_idle,
  Mmap2Stream_11___n__q0,
  Mmap2Stream_11___rmem11__q0,
  Mmap2Stream_11__ap_start,
  Mmap2Stream_11__ap_ready,
  Mmap2Stream_11__ap_done,
  Mmap2Stream_11__ap_idle,
  Mmap2Stream_12___n__q0,
  Mmap2Stream_12___rmem12__q0,
  Mmap2Stream_12__ap_start,
  Mmap2Stream_12__ap_ready,
  Mmap2Stream_12__ap_done,
  Mmap2Stream_12__ap_idle,
  Mmap2Stream_13___n__q0,
  Mmap2Stream_13___rmem13__q0,
  Mmap2Stream_13__ap_start,
  Mmap2Stream_13__ap_ready,
  Mmap2Stream_13__ap_done,
  Mmap2Stream_13__ap_idle,
  Mmap2Stream_14___n__q0,
  Mmap2Stream_14___rmem14__q0,
  Mmap2Stream_14__ap_start,
  Mmap2Stream_14__ap_ready,
  Mmap2Stream_14__ap_done,
  Mmap2Stream_14__ap_idle,
  Mmap2Stream_15___n__q0,
  Mmap2Stream_15___rmem15__q0,
  Mmap2Stream_15__ap_start,
  Mmap2Stream_15__ap_ready,
  Mmap2Stream_15__ap_done,
  Mmap2Stream_15__ap_idle,
  Mmap2Stream_16___n__q0,
  Mmap2Stream_16___rmem16__q0,
  Mmap2Stream_16__ap_start,
  Mmap2Stream_16__ap_ready,
  Mmap2Stream_16__ap_done,
  Mmap2Stream_16__ap_idle,
  Mmap2Stream_17___n__q0,
  Mmap2Stream_17___rmem17__q0,
  Mmap2Stream_17__ap_start,
  Mmap2Stream_17__ap_ready,
  Mmap2Stream_17__ap_done,
  Mmap2Stream_17__ap_idle,
  Mmap2Stream_18___n__q0,
  Mmap2Stream_18___rmem18__q0,
  Mmap2Stream_18__ap_start,
  Mmap2Stream_18__ap_ready,
  Mmap2Stream_18__ap_done,
  Mmap2Stream_18__ap_idle,
  Mmap2Stream_19___n__q0,
  Mmap2Stream_19___rmem19__q0,
  Mmap2Stream_19__ap_start,
  Mmap2Stream_19__ap_ready,
  Mmap2Stream_19__ap_done,
  Mmap2Stream_19__ap_idle,
  Mmap2Stream_20___n__q0,
  Mmap2Stream_20___rmem20__q0,
  Mmap2Stream_20__ap_start,
  Mmap2Stream_20__ap_ready,
  Mmap2Stream_20__ap_done,
  Mmap2Stream_20__ap_idle,
  Mmap2Stream_21___n__q0,
  Mmap2Stream_21___rmem21__q0,
  Mmap2Stream_21__ap_start,
  Mmap2Stream_21__ap_ready,
  Mmap2Stream_21__ap_done,
  Mmap2Stream_21__ap_idle,
  Mmap2Stream_22___n__q0,
  Mmap2Stream_22___rmem22__q0,
  Mmap2Stream_22__ap_start,
  Mmap2Stream_22__ap_ready,
  Mmap2Stream_22__ap_done,
  Mmap2Stream_22__ap_idle,
  Mmap2Stream_23___n__q0,
  Mmap2Stream_23___rmem23__q0,
  Mmap2Stream_23__ap_start,
  Mmap2Stream_23__ap_ready,
  Mmap2Stream_23__ap_done,
  Mmap2Stream_23__ap_idle,
  Mmap2Stream_24___n__q0,
  Mmap2Stream_24___rmem24__q0,
  Mmap2Stream_24__ap_start,
  Mmap2Stream_24__ap_ready,
  Mmap2Stream_24__ap_done,
  Mmap2Stream_24__ap_idle,
  Mmap2Stream_25___n__q0,
  Mmap2Stream_25___rmem25__q0,
  Mmap2Stream_25__ap_start,
  Mmap2Stream_25__ap_ready,
  Mmap2Stream_25__ap_done,
  Mmap2Stream_25__ap_idle,
  Mmap2Stream_26___n__q0,
  Mmap2Stream_26___rmem26__q0,
  Mmap2Stream_26__ap_start,
  Mmap2Stream_26__ap_ready,
  Mmap2Stream_26__ap_done,
  Mmap2Stream_26__ap_idle,
  Mmap2Stream_27___n__q0,
  Mmap2Stream_27___rmem27__q0,
  Mmap2Stream_27__ap_start,
  Mmap2Stream_27__ap_ready,
  Mmap2Stream_27__ap_done,
  Mmap2Stream_27__ap_idle,
  Mmap2Stream_28___n__q0,
  Mmap2Stream_28___rmem28__q0,
  Mmap2Stream_28__ap_start,
  Mmap2Stream_28__ap_ready,
  Mmap2Stream_28__ap_done,
  Mmap2Stream_28__ap_idle,
  Mmap2Stream_29___n__q0,
  Mmap2Stream_29___rmem29__q0,
  Mmap2Stream_29__ap_start,
  Mmap2Stream_29__ap_ready,
  Mmap2Stream_29__ap_done,
  Mmap2Stream_29__ap_idle,
  Stream2Mmap_0___n__q0,
  Stream2Mmap_0___wmem0__q0,
  Stream2Mmap_0__ap_start,
  Stream2Mmap_0__ap_ready,
  Stream2Mmap_0__ap_done,
  Stream2Mmap_0__ap_idle,
  yxor_0___n__q0,
  yxor_0__ap_start,
  yxor_0__ap_ready,
  yxor_0__ap_done,
  yxor_0__ap_idle,
  yxor_1___n__q0,
  yxor_1__ap_start,
  yxor_1__ap_ready,
  yxor_1__ap_done,
  yxor_1__ap_idle,
  yxor_2___n__q0,
  yxor_2__ap_start,
  yxor_2__ap_ready,
  yxor_2__ap_done,
  yxor_2__ap_idle,
  yxor_3___n__q0,
  yxor_3__ap_start,
  yxor_3__ap_ready,
  yxor_3__ap_done,
  yxor_3__ap_idle,
  yxor_4___n__q0,
  yxor_4__ap_start,
  yxor_4__ap_ready,
  yxor_4__ap_done,
  yxor_4__ap_idle,
  yxor_5___n__q0,
  yxor_5__ap_start,
  yxor_5__ap_ready,
  yxor_5__ap_done,
  yxor_5__ap_idle,
  yxor_6___n__q0,
  yxor_6__ap_start,
  yxor_6__ap_ready,
  yxor_6__ap_done,
  yxor_6__ap_idle,
  yxor_7___n__q0,
  yxor_7__ap_start,
  yxor_7__ap_ready,
  yxor_7__ap_done,
  yxor_7__ap_idle,
  yxor_8___n__q0,
  yxor_8__ap_start,
  yxor_8__ap_ready,
  yxor_8__ap_done,
  yxor_8__ap_idle,
  yxor_9___n__q0,
  yxor_9__ap_start,
  yxor_9__ap_ready,
  yxor_9__ap_done,
  yxor_9__ap_idle,
  yxor_10___n__q0,
  yxor_10__ap_start,
  yxor_10__ap_ready,
  yxor_10__ap_done,
  yxor_10__ap_idle,
  yxor_11___n__q0,
  yxor_11__ap_start,
  yxor_11__ap_ready,
  yxor_11__ap_done,
  yxor_11__ap_idle,
  yxor_12___n__q0,
  yxor_12__ap_start,
  yxor_12__ap_ready,
  yxor_12__ap_done,
  yxor_12__ap_idle,
  yxor_13___n__q0,
  yxor_13__ap_start,
  yxor_13__ap_ready,
  yxor_13__ap_done,
  yxor_13__ap_idle,
  yxor_14___n__q0,
  yxor_14__ap_start,
  yxor_14__ap_ready,
  yxor_14__ap_done,
  yxor_14__ap_idle,
  yxor_15___n__q0,
  yxor_15__ap_start,
  yxor_15__ap_ready,
  yxor_15__ap_done,
  yxor_15__ap_idle,
  yxor_16___n__q0,
  yxor_16__ap_start,
  yxor_16__ap_ready,
  yxor_16__ap_done,
  yxor_16__ap_idle,
  yxor_17___n__q0,
  yxor_17__ap_start,
  yxor_17__ap_ready,
  yxor_17__ap_done,
  yxor_17__ap_idle,
  yxor_18___n__q0,
  yxor_18__ap_start,
  yxor_18__ap_ready,
  yxor_18__ap_done,
  yxor_18__ap_idle,
  yxor_19___n__q0,
  yxor_19__ap_start,
  yxor_19__ap_ready,
  yxor_19__ap_done,
  yxor_19__ap_idle,
  yxor_20___n__q0,
  yxor_20__ap_start,
  yxor_20__ap_ready,
  yxor_20__ap_done,
  yxor_20__ap_idle,
  yxor_21___n__q0,
  yxor_21__ap_start,
  yxor_21__ap_ready,
  yxor_21__ap_done,
  yxor_21__ap_idle,
  yxor_22___n__q0,
  yxor_22__ap_start,
  yxor_22__ap_ready,
  yxor_22__ap_done,
  yxor_22__ap_idle,
  yxor_23___n__q0,
  yxor_23__ap_start,
  yxor_23__ap_ready,
  yxor_23__ap_done,
  yxor_23__ap_idle,
  yxor_24___n__q0,
  yxor_24__ap_start,
  yxor_24__ap_ready,
  yxor_24__ap_done,
  yxor_24__ap_idle,
  yxor_25___n__q0,
  yxor_25__ap_start,
  yxor_25__ap_ready,
  yxor_25__ap_done,
  yxor_25__ap_idle,
  yxor_26___n__q0,
  yxor_26__ap_start,
  yxor_26__ap_ready,
  yxor_26__ap_done,
  yxor_26__ap_idle,
  yxor_27___n__q0,
  yxor_27__ap_start,
  yxor_27__ap_ready,
  yxor_27__ap_done,
  yxor_27__ap_idle,
  yxor_28___n__q0,
  yxor_28__ap_start,
  yxor_28__ap_ready,
  yxor_28__ap_done,
  yxor_28__ap_idle
);

  // pragma RS clk port=ap_clk
  // pragma RS rst port=ap_rst_n active=low
  // pragma RS ap-ctrl ap_start=ap_start ap_done=ap_done ap_idle=ap_idle ap_ready=ap_ready scalar=(rmem0|rmem1|rmem2|rmem3|rmem4|rmem5|rmem6|rmem7|rmem8|rmem9|rmem10|rmem11|rmem12|rmem13|rmem14|rmem15|rmem16|rmem17|rmem18|rmem19|rmem20|rmem21|rmem22|rmem23|rmem24|rmem25|rmem26|rmem27|rmem28|rmem29|wmem0|n)
  // pragma RS ap-ctrl ap_start=Mmap2Stream_0__ap_start ap_done=Mmap2Stream_0__ap_done ap_idle=Mmap2Stream_0__ap_idle ap_ready=Mmap2Stream_0__ap_ready scalar=Mmap2Stream_0___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_1__ap_start ap_done=Mmap2Stream_1__ap_done ap_idle=Mmap2Stream_1__ap_idle ap_ready=Mmap2Stream_1__ap_ready scalar=Mmap2Stream_1___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_2__ap_start ap_done=Mmap2Stream_2__ap_done ap_idle=Mmap2Stream_2__ap_idle ap_ready=Mmap2Stream_2__ap_ready scalar=Mmap2Stream_2___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_3__ap_start ap_done=Mmap2Stream_3__ap_done ap_idle=Mmap2Stream_3__ap_idle ap_ready=Mmap2Stream_3__ap_ready scalar=Mmap2Stream_3___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_4__ap_start ap_done=Mmap2Stream_4__ap_done ap_idle=Mmap2Stream_4__ap_idle ap_ready=Mmap2Stream_4__ap_ready scalar=Mmap2Stream_4___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_5__ap_start ap_done=Mmap2Stream_5__ap_done ap_idle=Mmap2Stream_5__ap_idle ap_ready=Mmap2Stream_5__ap_ready scalar=Mmap2Stream_5___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_6__ap_start ap_done=Mmap2Stream_6__ap_done ap_idle=Mmap2Stream_6__ap_idle ap_ready=Mmap2Stream_6__ap_ready scalar=Mmap2Stream_6___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_7__ap_start ap_done=Mmap2Stream_7__ap_done ap_idle=Mmap2Stream_7__ap_idle ap_ready=Mmap2Stream_7__ap_ready scalar=Mmap2Stream_7___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_8__ap_start ap_done=Mmap2Stream_8__ap_done ap_idle=Mmap2Stream_8__ap_idle ap_ready=Mmap2Stream_8__ap_ready scalar=Mmap2Stream_8___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_9__ap_start ap_done=Mmap2Stream_9__ap_done ap_idle=Mmap2Stream_9__ap_idle ap_ready=Mmap2Stream_9__ap_ready scalar=Mmap2Stream_9___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_10__ap_start ap_done=Mmap2Stream_10__ap_done ap_idle=Mmap2Stream_10__ap_idle ap_ready=Mmap2Stream_10__ap_ready scalar=Mmap2Stream_10___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_11__ap_start ap_done=Mmap2Stream_11__ap_done ap_idle=Mmap2Stream_11__ap_idle ap_ready=Mmap2Stream_11__ap_ready scalar=Mmap2Stream_11___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_12__ap_start ap_done=Mmap2Stream_12__ap_done ap_idle=Mmap2Stream_12__ap_idle ap_ready=Mmap2Stream_12__ap_ready scalar=Mmap2Stream_12___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_13__ap_start ap_done=Mmap2Stream_13__ap_done ap_idle=Mmap2Stream_13__ap_idle ap_ready=Mmap2Stream_13__ap_ready scalar=Mmap2Stream_13___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_14__ap_start ap_done=Mmap2Stream_14__ap_done ap_idle=Mmap2Stream_14__ap_idle ap_ready=Mmap2Stream_14__ap_ready scalar=Mmap2Stream_14___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_15__ap_start ap_done=Mmap2Stream_15__ap_done ap_idle=Mmap2Stream_15__ap_idle ap_ready=Mmap2Stream_15__ap_ready scalar=Mmap2Stream_15___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_16__ap_start ap_done=Mmap2Stream_16__ap_done ap_idle=Mmap2Stream_16__ap_idle ap_ready=Mmap2Stream_16__ap_ready scalar=Mmap2Stream_16___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_17__ap_start ap_done=Mmap2Stream_17__ap_done ap_idle=Mmap2Stream_17__ap_idle ap_ready=Mmap2Stream_17__ap_ready scalar=Mmap2Stream_17___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_18__ap_start ap_done=Mmap2Stream_18__ap_done ap_idle=Mmap2Stream_18__ap_idle ap_ready=Mmap2Stream_18__ap_ready scalar=Mmap2Stream_18___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_19__ap_start ap_done=Mmap2Stream_19__ap_done ap_idle=Mmap2Stream_19__ap_idle ap_ready=Mmap2Stream_19__ap_ready scalar=Mmap2Stream_19___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_20__ap_start ap_done=Mmap2Stream_20__ap_done ap_idle=Mmap2Stream_20__ap_idle ap_ready=Mmap2Stream_20__ap_ready scalar=Mmap2Stream_20___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_21__ap_start ap_done=Mmap2Stream_21__ap_done ap_idle=Mmap2Stream_21__ap_idle ap_ready=Mmap2Stream_21__ap_ready scalar=Mmap2Stream_21___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_22__ap_start ap_done=Mmap2Stream_22__ap_done ap_idle=Mmap2Stream_22__ap_idle ap_ready=Mmap2Stream_22__ap_ready scalar=Mmap2Stream_22___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_23__ap_start ap_done=Mmap2Stream_23__ap_done ap_idle=Mmap2Stream_23__ap_idle ap_ready=Mmap2Stream_23__ap_ready scalar=Mmap2Stream_23___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_24__ap_start ap_done=Mmap2Stream_24__ap_done ap_idle=Mmap2Stream_24__ap_idle ap_ready=Mmap2Stream_24__ap_ready scalar=Mmap2Stream_24___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_25__ap_start ap_done=Mmap2Stream_25__ap_done ap_idle=Mmap2Stream_25__ap_idle ap_ready=Mmap2Stream_25__ap_ready scalar=Mmap2Stream_25___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_26__ap_start ap_done=Mmap2Stream_26__ap_done ap_idle=Mmap2Stream_26__ap_idle ap_ready=Mmap2Stream_26__ap_ready scalar=Mmap2Stream_26___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_27__ap_start ap_done=Mmap2Stream_27__ap_done ap_idle=Mmap2Stream_27__ap_idle ap_ready=Mmap2Stream_27__ap_ready scalar=Mmap2Stream_27___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_28__ap_start ap_done=Mmap2Stream_28__ap_done ap_idle=Mmap2Stream_28__ap_idle ap_ready=Mmap2Stream_28__ap_ready scalar=Mmap2Stream_28___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_29__ap_start ap_done=Mmap2Stream_29__ap_done ap_idle=Mmap2Stream_29__ap_idle ap_ready=Mmap2Stream_29__ap_ready scalar=Mmap2Stream_29___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_0__ap_start ap_done=Stream2Mmap_0__ap_done ap_idle=Stream2Mmap_0__ap_idle ap_ready=Stream2Mmap_0__ap_ready scalar=Stream2Mmap_0___.*
  // pragma RS ap-ctrl ap_start=yxor_0__ap_start ap_done=yxor_0__ap_done ap_idle=yxor_0__ap_idle ap_ready=yxor_0__ap_ready scalar=yxor_0___.*
  // pragma RS ap-ctrl ap_start=yxor_1__ap_start ap_done=yxor_1__ap_done ap_idle=yxor_1__ap_idle ap_ready=yxor_1__ap_ready scalar=yxor_1___.*
  // pragma RS ap-ctrl ap_start=yxor_2__ap_start ap_done=yxor_2__ap_done ap_idle=yxor_2__ap_idle ap_ready=yxor_2__ap_ready scalar=yxor_2___.*
  // pragma RS ap-ctrl ap_start=yxor_3__ap_start ap_done=yxor_3__ap_done ap_idle=yxor_3__ap_idle ap_ready=yxor_3__ap_ready scalar=yxor_3___.*
  // pragma RS ap-ctrl ap_start=yxor_4__ap_start ap_done=yxor_4__ap_done ap_idle=yxor_4__ap_idle ap_ready=yxor_4__ap_ready scalar=yxor_4___.*
  // pragma RS ap-ctrl ap_start=yxor_5__ap_start ap_done=yxor_5__ap_done ap_idle=yxor_5__ap_idle ap_ready=yxor_5__ap_ready scalar=yxor_5___.*
  // pragma RS ap-ctrl ap_start=yxor_6__ap_start ap_done=yxor_6__ap_done ap_idle=yxor_6__ap_idle ap_ready=yxor_6__ap_ready scalar=yxor_6___.*
  // pragma RS ap-ctrl ap_start=yxor_7__ap_start ap_done=yxor_7__ap_done ap_idle=yxor_7__ap_idle ap_ready=yxor_7__ap_ready scalar=yxor_7___.*
  // pragma RS ap-ctrl ap_start=yxor_8__ap_start ap_done=yxor_8__ap_done ap_idle=yxor_8__ap_idle ap_ready=yxor_8__ap_ready scalar=yxor_8___.*
  // pragma RS ap-ctrl ap_start=yxor_9__ap_start ap_done=yxor_9__ap_done ap_idle=yxor_9__ap_idle ap_ready=yxor_9__ap_ready scalar=yxor_9___.*
  // pragma RS ap-ctrl ap_start=yxor_10__ap_start ap_done=yxor_10__ap_done ap_idle=yxor_10__ap_idle ap_ready=yxor_10__ap_ready scalar=yxor_10___.*
  // pragma RS ap-ctrl ap_start=yxor_11__ap_start ap_done=yxor_11__ap_done ap_idle=yxor_11__ap_idle ap_ready=yxor_11__ap_ready scalar=yxor_11___.*
  // pragma RS ap-ctrl ap_start=yxor_12__ap_start ap_done=yxor_12__ap_done ap_idle=yxor_12__ap_idle ap_ready=yxor_12__ap_ready scalar=yxor_12___.*
  // pragma RS ap-ctrl ap_start=yxor_13__ap_start ap_done=yxor_13__ap_done ap_idle=yxor_13__ap_idle ap_ready=yxor_13__ap_ready scalar=yxor_13___.*
  // pragma RS ap-ctrl ap_start=yxor_14__ap_start ap_done=yxor_14__ap_done ap_idle=yxor_14__ap_idle ap_ready=yxor_14__ap_ready scalar=yxor_14___.*
  // pragma RS ap-ctrl ap_start=yxor_15__ap_start ap_done=yxor_15__ap_done ap_idle=yxor_15__ap_idle ap_ready=yxor_15__ap_ready scalar=yxor_15___.*
  // pragma RS ap-ctrl ap_start=yxor_16__ap_start ap_done=yxor_16__ap_done ap_idle=yxor_16__ap_idle ap_ready=yxor_16__ap_ready scalar=yxor_16___.*
  // pragma RS ap-ctrl ap_start=yxor_17__ap_start ap_done=yxor_17__ap_done ap_idle=yxor_17__ap_idle ap_ready=yxor_17__ap_ready scalar=yxor_17___.*
  // pragma RS ap-ctrl ap_start=yxor_18__ap_start ap_done=yxor_18__ap_done ap_idle=yxor_18__ap_idle ap_ready=yxor_18__ap_ready scalar=yxor_18___.*
  // pragma RS ap-ctrl ap_start=yxor_19__ap_start ap_done=yxor_19__ap_done ap_idle=yxor_19__ap_idle ap_ready=yxor_19__ap_ready scalar=yxor_19___.*
  // pragma RS ap-ctrl ap_start=yxor_20__ap_start ap_done=yxor_20__ap_done ap_idle=yxor_20__ap_idle ap_ready=yxor_20__ap_ready scalar=yxor_20___.*
  // pragma RS ap-ctrl ap_start=yxor_21__ap_start ap_done=yxor_21__ap_done ap_idle=yxor_21__ap_idle ap_ready=yxor_21__ap_ready scalar=yxor_21___.*
  // pragma RS ap-ctrl ap_start=yxor_22__ap_start ap_done=yxor_22__ap_done ap_idle=yxor_22__ap_idle ap_ready=yxor_22__ap_ready scalar=yxor_22___.*
  // pragma RS ap-ctrl ap_start=yxor_23__ap_start ap_done=yxor_23__ap_done ap_idle=yxor_23__ap_idle ap_ready=yxor_23__ap_ready scalar=yxor_23___.*
  // pragma RS ap-ctrl ap_start=yxor_24__ap_start ap_done=yxor_24__ap_done ap_idle=yxor_24__ap_idle ap_ready=yxor_24__ap_ready scalar=yxor_24___.*
  // pragma RS ap-ctrl ap_start=yxor_25__ap_start ap_done=yxor_25__ap_done ap_idle=yxor_25__ap_idle ap_ready=yxor_25__ap_ready scalar=yxor_25___.*
  // pragma RS ap-ctrl ap_start=yxor_26__ap_start ap_done=yxor_26__ap_done ap_idle=yxor_26__ap_idle ap_ready=yxor_26__ap_ready scalar=yxor_26___.*
  // pragma RS ap-ctrl ap_start=yxor_27__ap_start ap_done=yxor_27__ap_done ap_idle=yxor_27__ap_idle ap_ready=yxor_27__ap_ready scalar=yxor_27___.*
  // pragma RS ap-ctrl ap_start=yxor_28__ap_start ap_done=yxor_28__ap_done ap_idle=yxor_28__ap_idle ap_ready=yxor_28__ap_ready scalar=yxor_28___.*

  input ap_clk;
  input ap_rst_n;
  input ap_start;
  output ap_ready;
  output ap_done;
  output ap_idle;
  input [63:0] n;
  input [63:0] rmem0;
  input [63:0] rmem1;
  input [63:0] rmem2;
  input [63:0] rmem3;
  input [63:0] rmem4;
  input [63:0] rmem5;
  input [63:0] rmem6;
  input [63:0] rmem7;
  input [63:0] rmem8;
  input [63:0] rmem9;
  input [63:0] rmem10;
  input [63:0] rmem11;
  input [63:0] rmem12;
  input [63:0] rmem13;
  input [63:0] rmem14;
  input [63:0] rmem15;
  input [63:0] rmem16;
  input [63:0] rmem17;
  input [63:0] rmem18;
  input [63:0] rmem19;
  input [63:0] rmem20;
  input [63:0] rmem21;
  input [63:0] rmem22;
  input [63:0] rmem23;
  input [63:0] rmem24;
  input [63:0] rmem25;
  input [63:0] rmem26;
  input [63:0] rmem27;
  input [63:0] rmem28;
  input [63:0] rmem29;
  input [63:0] wmem0;
  output [63:0] Mmap2Stream_0___n__q0;
  output [63:0] Mmap2Stream_0___rmem0__q0;
  output Mmap2Stream_0__ap_start;
  input Mmap2Stream_0__ap_ready;
  input Mmap2Stream_0__ap_done;
  input Mmap2Stream_0__ap_idle;
  output [63:0] Mmap2Stream_1___n__q0;
  output [63:0] Mmap2Stream_1___rmem1__q0;
  output Mmap2Stream_1__ap_start;
  input Mmap2Stream_1__ap_ready;
  input Mmap2Stream_1__ap_done;
  input Mmap2Stream_1__ap_idle;
  output [63:0] Mmap2Stream_2___n__q0;
  output [63:0] Mmap2Stream_2___rmem2__q0;
  output Mmap2Stream_2__ap_start;
  input Mmap2Stream_2__ap_ready;
  input Mmap2Stream_2__ap_done;
  input Mmap2Stream_2__ap_idle;
  output [63:0] Mmap2Stream_3___n__q0;
  output [63:0] Mmap2Stream_3___rmem3__q0;
  output Mmap2Stream_3__ap_start;
  input Mmap2Stream_3__ap_ready;
  input Mmap2Stream_3__ap_done;
  input Mmap2Stream_3__ap_idle;
  output [63:0] Mmap2Stream_4___n__q0;
  output [63:0] Mmap2Stream_4___rmem4__q0;
  output Mmap2Stream_4__ap_start;
  input Mmap2Stream_4__ap_ready;
  input Mmap2Stream_4__ap_done;
  input Mmap2Stream_4__ap_idle;
  output [63:0] Mmap2Stream_5___n__q0;
  output [63:0] Mmap2Stream_5___rmem5__q0;
  output Mmap2Stream_5__ap_start;
  input Mmap2Stream_5__ap_ready;
  input Mmap2Stream_5__ap_done;
  input Mmap2Stream_5__ap_idle;
  output [63:0] Mmap2Stream_6___n__q0;
  output [63:0] Mmap2Stream_6___rmem6__q0;
  output Mmap2Stream_6__ap_start;
  input Mmap2Stream_6__ap_ready;
  input Mmap2Stream_6__ap_done;
  input Mmap2Stream_6__ap_idle;
  output [63:0] Mmap2Stream_7___n__q0;
  output [63:0] Mmap2Stream_7___rmem7__q0;
  output Mmap2Stream_7__ap_start;
  input Mmap2Stream_7__ap_ready;
  input Mmap2Stream_7__ap_done;
  input Mmap2Stream_7__ap_idle;
  output [63:0] Mmap2Stream_8___n__q0;
  output [63:0] Mmap2Stream_8___rmem8__q0;
  output Mmap2Stream_8__ap_start;
  input Mmap2Stream_8__ap_ready;
  input Mmap2Stream_8__ap_done;
  input Mmap2Stream_8__ap_idle;
  output [63:0] Mmap2Stream_9___n__q0;
  output [63:0] Mmap2Stream_9___rmem9__q0;
  output Mmap2Stream_9__ap_start;
  input Mmap2Stream_9__ap_ready;
  input Mmap2Stream_9__ap_done;
  input Mmap2Stream_9__ap_idle;
  output [63:0] Mmap2Stream_10___n__q0;
  output [63:0] Mmap2Stream_10___rmem10__q0;
  output Mmap2Stream_10__ap_start;
  input Mmap2Stream_10__ap_ready;
  input Mmap2Stream_10__ap_done;
  input Mmap2Stream_10__ap_idle;
  output [63:0] Mmap2Stream_11___n__q0;
  output [63:0] Mmap2Stream_11___rmem11__q0;
  output Mmap2Stream_11__ap_start;
  input Mmap2Stream_11__ap_ready;
  input Mmap2Stream_11__ap_done;
  input Mmap2Stream_11__ap_idle;
  output [63:0] Mmap2Stream_12___n__q0;
  output [63:0] Mmap2Stream_12___rmem12__q0;
  output Mmap2Stream_12__ap_start;
  input Mmap2Stream_12__ap_ready;
  input Mmap2Stream_12__ap_done;
  input Mmap2Stream_12__ap_idle;
  output [63:0] Mmap2Stream_13___n__q0;
  output [63:0] Mmap2Stream_13___rmem13__q0;
  output Mmap2Stream_13__ap_start;
  input Mmap2Stream_13__ap_ready;
  input Mmap2Stream_13__ap_done;
  input Mmap2Stream_13__ap_idle;
  output [63:0] Mmap2Stream_14___n__q0;
  output [63:0] Mmap2Stream_14___rmem14__q0;
  output Mmap2Stream_14__ap_start;
  input Mmap2Stream_14__ap_ready;
  input Mmap2Stream_14__ap_done;
  input Mmap2Stream_14__ap_idle;
  output [63:0] Mmap2Stream_15___n__q0;
  output [63:0] Mmap2Stream_15___rmem15__q0;
  output Mmap2Stream_15__ap_start;
  input Mmap2Stream_15__ap_ready;
  input Mmap2Stream_15__ap_done;
  input Mmap2Stream_15__ap_idle;
  output [63:0] Mmap2Stream_16___n__q0;
  output [63:0] Mmap2Stream_16___rmem16__q0;
  output Mmap2Stream_16__ap_start;
  input Mmap2Stream_16__ap_ready;
  input Mmap2Stream_16__ap_done;
  input Mmap2Stream_16__ap_idle;
  output [63:0] Mmap2Stream_17___n__q0;
  output [63:0] Mmap2Stream_17___rmem17__q0;
  output Mmap2Stream_17__ap_start;
  input Mmap2Stream_17__ap_ready;
  input Mmap2Stream_17__ap_done;
  input Mmap2Stream_17__ap_idle;
  output [63:0] Mmap2Stream_18___n__q0;
  output [63:0] Mmap2Stream_18___rmem18__q0;
  output Mmap2Stream_18__ap_start;
  input Mmap2Stream_18__ap_ready;
  input Mmap2Stream_18__ap_done;
  input Mmap2Stream_18__ap_idle;
  output [63:0] Mmap2Stream_19___n__q0;
  output [63:0] Mmap2Stream_19___rmem19__q0;
  output Mmap2Stream_19__ap_start;
  input Mmap2Stream_19__ap_ready;
  input Mmap2Stream_19__ap_done;
  input Mmap2Stream_19__ap_idle;
  output [63:0] Mmap2Stream_20___n__q0;
  output [63:0] Mmap2Stream_20___rmem20__q0;
  output Mmap2Stream_20__ap_start;
  input Mmap2Stream_20__ap_ready;
  input Mmap2Stream_20__ap_done;
  input Mmap2Stream_20__ap_idle;
  output [63:0] Mmap2Stream_21___n__q0;
  output [63:0] Mmap2Stream_21___rmem21__q0;
  output Mmap2Stream_21__ap_start;
  input Mmap2Stream_21__ap_ready;
  input Mmap2Stream_21__ap_done;
  input Mmap2Stream_21__ap_idle;
  output [63:0] Mmap2Stream_22___n__q0;
  output [63:0] Mmap2Stream_22___rmem22__q0;
  output Mmap2Stream_22__ap_start;
  input Mmap2Stream_22__ap_ready;
  input Mmap2Stream_22__ap_done;
  input Mmap2Stream_22__ap_idle;
  output [63:0] Mmap2Stream_23___n__q0;
  output [63:0] Mmap2Stream_23___rmem23__q0;
  output Mmap2Stream_23__ap_start;
  input Mmap2Stream_23__ap_ready;
  input Mmap2Stream_23__ap_done;
  input Mmap2Stream_23__ap_idle;
  output [63:0] Mmap2Stream_24___n__q0;
  output [63:0] Mmap2Stream_24___rmem24__q0;
  output Mmap2Stream_24__ap_start;
  input Mmap2Stream_24__ap_ready;
  input Mmap2Stream_24__ap_done;
  input Mmap2Stream_24__ap_idle;
  output [63:0] Mmap2Stream_25___n__q0;
  output [63:0] Mmap2Stream_25___rmem25__q0;
  output Mmap2Stream_25__ap_start;
  input Mmap2Stream_25__ap_ready;
  input Mmap2Stream_25__ap_done;
  input Mmap2Stream_25__ap_idle;
  output [63:0] Mmap2Stream_26___n__q0;
  output [63:0] Mmap2Stream_26___rmem26__q0;
  output Mmap2Stream_26__ap_start;
  input Mmap2Stream_26__ap_ready;
  input Mmap2Stream_26__ap_done;
  input Mmap2Stream_26__ap_idle;
  output [63:0] Mmap2Stream_27___n__q0;
  output [63:0] Mmap2Stream_27___rmem27__q0;
  output Mmap2Stream_27__ap_start;
  input Mmap2Stream_27__ap_ready;
  input Mmap2Stream_27__ap_done;
  input Mmap2Stream_27__ap_idle;
  output [63:0] Mmap2Stream_28___n__q0;
  output [63:0] Mmap2Stream_28___rmem28__q0;
  output Mmap2Stream_28__ap_start;
  input Mmap2Stream_28__ap_ready;
  input Mmap2Stream_28__ap_done;
  input Mmap2Stream_28__ap_idle;
  output [63:0] Mmap2Stream_29___n__q0;
  output [63:0] Mmap2Stream_29___rmem29__q0;
  output Mmap2Stream_29__ap_start;
  input Mmap2Stream_29__ap_ready;
  input Mmap2Stream_29__ap_done;
  input Mmap2Stream_29__ap_idle;
  output [63:0] Stream2Mmap_0___n__q0;
  output [63:0] Stream2Mmap_0___wmem0__q0;
  output Stream2Mmap_0__ap_start;
  input Stream2Mmap_0__ap_ready;
  input Stream2Mmap_0__ap_done;
  input Stream2Mmap_0__ap_idle;
  output [63:0] yxor_0___n__q0;
  output yxor_0__ap_start;
  input yxor_0__ap_ready;
  input yxor_0__ap_done;
  input yxor_0__ap_idle;
  output [63:0] yxor_1___n__q0;
  output yxor_1__ap_start;
  input yxor_1__ap_ready;
  input yxor_1__ap_done;
  input yxor_1__ap_idle;
  output [63:0] yxor_2___n__q0;
  output yxor_2__ap_start;
  input yxor_2__ap_ready;
  input yxor_2__ap_done;
  input yxor_2__ap_idle;
  output [63:0] yxor_3___n__q0;
  output yxor_3__ap_start;
  input yxor_3__ap_ready;
  input yxor_3__ap_done;
  input yxor_3__ap_idle;
  output [63:0] yxor_4___n__q0;
  output yxor_4__ap_start;
  input yxor_4__ap_ready;
  input yxor_4__ap_done;
  input yxor_4__ap_idle;
  output [63:0] yxor_5___n__q0;
  output yxor_5__ap_start;
  input yxor_5__ap_ready;
  input yxor_5__ap_done;
  input yxor_5__ap_idle;
  output [63:0] yxor_6___n__q0;
  output yxor_6__ap_start;
  input yxor_6__ap_ready;
  input yxor_6__ap_done;
  input yxor_6__ap_idle;
  output [63:0] yxor_7___n__q0;
  output yxor_7__ap_start;
  input yxor_7__ap_ready;
  input yxor_7__ap_done;
  input yxor_7__ap_idle;
  output [63:0] yxor_8___n__q0;
  output yxor_8__ap_start;
  input yxor_8__ap_ready;
  input yxor_8__ap_done;
  input yxor_8__ap_idle;
  output [63:0] yxor_9___n__q0;
  output yxor_9__ap_start;
  input yxor_9__ap_ready;
  input yxor_9__ap_done;
  input yxor_9__ap_idle;
  output [63:0] yxor_10___n__q0;
  output yxor_10__ap_start;
  input yxor_10__ap_ready;
  input yxor_10__ap_done;
  input yxor_10__ap_idle;
  output [63:0] yxor_11___n__q0;
  output yxor_11__ap_start;
  input yxor_11__ap_ready;
  input yxor_11__ap_done;
  input yxor_11__ap_idle;
  output [63:0] yxor_12___n__q0;
  output yxor_12__ap_start;
  input yxor_12__ap_ready;
  input yxor_12__ap_done;
  input yxor_12__ap_idle;
  output [63:0] yxor_13___n__q0;
  output yxor_13__ap_start;
  input yxor_13__ap_ready;
  input yxor_13__ap_done;
  input yxor_13__ap_idle;
  output [63:0] yxor_14___n__q0;
  output yxor_14__ap_start;
  input yxor_14__ap_ready;
  input yxor_14__ap_done;
  input yxor_14__ap_idle;
  output [63:0] yxor_15___n__q0;
  output yxor_15__ap_start;
  input yxor_15__ap_ready;
  input yxor_15__ap_done;
  input yxor_15__ap_idle;
  output [63:0] yxor_16___n__q0;
  output yxor_16__ap_start;
  input yxor_16__ap_ready;
  input yxor_16__ap_done;
  input yxor_16__ap_idle;
  output [63:0] yxor_17___n__q0;
  output yxor_17__ap_start;
  input yxor_17__ap_ready;
  input yxor_17__ap_done;
  input yxor_17__ap_idle;
  output [63:0] yxor_18___n__q0;
  output yxor_18__ap_start;
  input yxor_18__ap_ready;
  input yxor_18__ap_done;
  input yxor_18__ap_idle;
  output [63:0] yxor_19___n__q0;
  output yxor_19__ap_start;
  input yxor_19__ap_ready;
  input yxor_19__ap_done;
  input yxor_19__ap_idle;
  output [63:0] yxor_20___n__q0;
  output yxor_20__ap_start;
  input yxor_20__ap_ready;
  input yxor_20__ap_done;
  input yxor_20__ap_idle;
  output [63:0] yxor_21___n__q0;
  output yxor_21__ap_start;
  input yxor_21__ap_ready;
  input yxor_21__ap_done;
  input yxor_21__ap_idle;
  output [63:0] yxor_22___n__q0;
  output yxor_22__ap_start;
  input yxor_22__ap_ready;
  input yxor_22__ap_done;
  input yxor_22__ap_idle;
  output [63:0] yxor_23___n__q0;
  output yxor_23__ap_start;
  input yxor_23__ap_ready;
  input yxor_23__ap_done;
  input yxor_23__ap_idle;
  output [63:0] yxor_24___n__q0;
  output yxor_24__ap_start;
  input yxor_24__ap_ready;
  input yxor_24__ap_done;
  input yxor_24__ap_idle;
  output [63:0] yxor_25___n__q0;
  output yxor_25__ap_start;
  input yxor_25__ap_ready;
  input yxor_25__ap_done;
  input yxor_25__ap_idle;
  output [63:0] yxor_26___n__q0;
  output yxor_26__ap_start;
  input yxor_26__ap_ready;
  input yxor_26__ap_done;
  input yxor_26__ap_idle;
  output [63:0] yxor_27___n__q0;
  output yxor_27__ap_start;
  input yxor_27__ap_ready;
  input yxor_27__ap_done;
  input yxor_27__ap_idle;
  output [63:0] yxor_28___n__q0;
  output yxor_28__ap_start;
  input yxor_28__ap_ready;
  input yxor_28__ap_done;
  input yxor_28__ap_idle;
  wire [63:0] Mmap2Stream_0___n__q0;
  wire [63:0] Mmap2Stream_0___rmem0__q0;
  wire Mmap2Stream_0__ap_start_global__q0;
  wire Mmap2Stream_0__is_done__q0;
  wire Mmap2Stream_0__ap_done_global__q0;
  wire Mmap2Stream_0__ap_start;
  wire Mmap2Stream_0__ap_ready;
  wire Mmap2Stream_0__ap_done;
  wire Mmap2Stream_0__ap_idle;
  reg [1:0] Mmap2Stream_0__state;
  wire [63:0] Mmap2Stream_1___n__q0;
  wire [63:0] Mmap2Stream_1___rmem1__q0;
  wire Mmap2Stream_1__ap_start_global__q0;
  wire Mmap2Stream_1__is_done__q0;
  wire Mmap2Stream_1__ap_done_global__q0;
  wire Mmap2Stream_1__ap_start;
  wire Mmap2Stream_1__ap_ready;
  wire Mmap2Stream_1__ap_done;
  wire Mmap2Stream_1__ap_idle;
  reg [1:0] Mmap2Stream_1__state;
  wire [63:0] Mmap2Stream_2___n__q0;
  wire [63:0] Mmap2Stream_2___rmem2__q0;
  wire Mmap2Stream_2__ap_start_global__q0;
  wire Mmap2Stream_2__is_done__q0;
  wire Mmap2Stream_2__ap_done_global__q0;
  wire Mmap2Stream_2__ap_start;
  wire Mmap2Stream_2__ap_ready;
  wire Mmap2Stream_2__ap_done;
  wire Mmap2Stream_2__ap_idle;
  reg [1:0] Mmap2Stream_2__state;
  wire [63:0] Mmap2Stream_3___n__q0;
  wire [63:0] Mmap2Stream_3___rmem3__q0;
  wire Mmap2Stream_3__ap_start_global__q0;
  wire Mmap2Stream_3__is_done__q0;
  wire Mmap2Stream_3__ap_done_global__q0;
  wire Mmap2Stream_3__ap_start;
  wire Mmap2Stream_3__ap_ready;
  wire Mmap2Stream_3__ap_done;
  wire Mmap2Stream_3__ap_idle;
  reg [1:0] Mmap2Stream_3__state;
  wire [63:0] Mmap2Stream_4___n__q0;
  wire [63:0] Mmap2Stream_4___rmem4__q0;
  wire Mmap2Stream_4__ap_start_global__q0;
  wire Mmap2Stream_4__is_done__q0;
  wire Mmap2Stream_4__ap_done_global__q0;
  wire Mmap2Stream_4__ap_start;
  wire Mmap2Stream_4__ap_ready;
  wire Mmap2Stream_4__ap_done;
  wire Mmap2Stream_4__ap_idle;
  reg [1:0] Mmap2Stream_4__state;
  wire [63:0] Mmap2Stream_5___n__q0;
  wire [63:0] Mmap2Stream_5___rmem5__q0;
  wire Mmap2Stream_5__ap_start_global__q0;
  wire Mmap2Stream_5__is_done__q0;
  wire Mmap2Stream_5__ap_done_global__q0;
  wire Mmap2Stream_5__ap_start;
  wire Mmap2Stream_5__ap_ready;
  wire Mmap2Stream_5__ap_done;
  wire Mmap2Stream_5__ap_idle;
  reg [1:0] Mmap2Stream_5__state;
  wire [63:0] Mmap2Stream_6___n__q0;
  wire [63:0] Mmap2Stream_6___rmem6__q0;
  wire Mmap2Stream_6__ap_start_global__q0;
  wire Mmap2Stream_6__is_done__q0;
  wire Mmap2Stream_6__ap_done_global__q0;
  wire Mmap2Stream_6__ap_start;
  wire Mmap2Stream_6__ap_ready;
  wire Mmap2Stream_6__ap_done;
  wire Mmap2Stream_6__ap_idle;
  reg [1:0] Mmap2Stream_6__state;
  wire [63:0] Mmap2Stream_7___n__q0;
  wire [63:0] Mmap2Stream_7___rmem7__q0;
  wire Mmap2Stream_7__ap_start_global__q0;
  wire Mmap2Stream_7__is_done__q0;
  wire Mmap2Stream_7__ap_done_global__q0;
  wire Mmap2Stream_7__ap_start;
  wire Mmap2Stream_7__ap_ready;
  wire Mmap2Stream_7__ap_done;
  wire Mmap2Stream_7__ap_idle;
  reg [1:0] Mmap2Stream_7__state;
  wire [63:0] Mmap2Stream_8___n__q0;
  wire [63:0] Mmap2Stream_8___rmem8__q0;
  wire Mmap2Stream_8__ap_start_global__q0;
  wire Mmap2Stream_8__is_done__q0;
  wire Mmap2Stream_8__ap_done_global__q0;
  wire Mmap2Stream_8__ap_start;
  wire Mmap2Stream_8__ap_ready;
  wire Mmap2Stream_8__ap_done;
  wire Mmap2Stream_8__ap_idle;
  reg [1:0] Mmap2Stream_8__state;
  wire [63:0] Mmap2Stream_9___n__q0;
  wire [63:0] Mmap2Stream_9___rmem9__q0;
  wire Mmap2Stream_9__ap_start_global__q0;
  wire Mmap2Stream_9__is_done__q0;
  wire Mmap2Stream_9__ap_done_global__q0;
  wire Mmap2Stream_9__ap_start;
  wire Mmap2Stream_9__ap_ready;
  wire Mmap2Stream_9__ap_done;
  wire Mmap2Stream_9__ap_idle;
  reg [1:0] Mmap2Stream_9__state;
  wire [63:0] Mmap2Stream_10___n__q0;
  wire [63:0] Mmap2Stream_10___rmem10__q0;
  wire Mmap2Stream_10__ap_start_global__q0;
  wire Mmap2Stream_10__is_done__q0;
  wire Mmap2Stream_10__ap_done_global__q0;
  wire Mmap2Stream_10__ap_start;
  wire Mmap2Stream_10__ap_ready;
  wire Mmap2Stream_10__ap_done;
  wire Mmap2Stream_10__ap_idle;
  reg [1:0] Mmap2Stream_10__state;
  wire [63:0] Mmap2Stream_11___n__q0;
  wire [63:0] Mmap2Stream_11___rmem11__q0;
  wire Mmap2Stream_11__ap_start_global__q0;
  wire Mmap2Stream_11__is_done__q0;
  wire Mmap2Stream_11__ap_done_global__q0;
  wire Mmap2Stream_11__ap_start;
  wire Mmap2Stream_11__ap_ready;
  wire Mmap2Stream_11__ap_done;
  wire Mmap2Stream_11__ap_idle;
  reg [1:0] Mmap2Stream_11__state;
  wire [63:0] Mmap2Stream_12___n__q0;
  wire [63:0] Mmap2Stream_12___rmem12__q0;
  wire Mmap2Stream_12__ap_start_global__q0;
  wire Mmap2Stream_12__is_done__q0;
  wire Mmap2Stream_12__ap_done_global__q0;
  wire Mmap2Stream_12__ap_start;
  wire Mmap2Stream_12__ap_ready;
  wire Mmap2Stream_12__ap_done;
  wire Mmap2Stream_12__ap_idle;
  reg [1:0] Mmap2Stream_12__state;
  wire [63:0] Mmap2Stream_13___n__q0;
  wire [63:0] Mmap2Stream_13___rmem13__q0;
  wire Mmap2Stream_13__ap_start_global__q0;
  wire Mmap2Stream_13__is_done__q0;
  wire Mmap2Stream_13__ap_done_global__q0;
  wire Mmap2Stream_13__ap_start;
  wire Mmap2Stream_13__ap_ready;
  wire Mmap2Stream_13__ap_done;
  wire Mmap2Stream_13__ap_idle;
  reg [1:0] Mmap2Stream_13__state;
  wire [63:0] Mmap2Stream_14___n__q0;
  wire [63:0] Mmap2Stream_14___rmem14__q0;
  wire Mmap2Stream_14__ap_start_global__q0;
  wire Mmap2Stream_14__is_done__q0;
  wire Mmap2Stream_14__ap_done_global__q0;
  wire Mmap2Stream_14__ap_start;
  wire Mmap2Stream_14__ap_ready;
  wire Mmap2Stream_14__ap_done;
  wire Mmap2Stream_14__ap_idle;
  reg [1:0] Mmap2Stream_14__state;
  wire [63:0] Mmap2Stream_15___n__q0;
  wire [63:0] Mmap2Stream_15___rmem15__q0;
  wire Mmap2Stream_15__ap_start_global__q0;
  wire Mmap2Stream_15__is_done__q0;
  wire Mmap2Stream_15__ap_done_global__q0;
  wire Mmap2Stream_15__ap_start;
  wire Mmap2Stream_15__ap_ready;
  wire Mmap2Stream_15__ap_done;
  wire Mmap2Stream_15__ap_idle;
  reg [1:0] Mmap2Stream_15__state;
  wire [63:0] Mmap2Stream_16___n__q0;
  wire [63:0] Mmap2Stream_16___rmem16__q0;
  wire Mmap2Stream_16__ap_start_global__q0;
  wire Mmap2Stream_16__is_done__q0;
  wire Mmap2Stream_16__ap_done_global__q0;
  wire Mmap2Stream_16__ap_start;
  wire Mmap2Stream_16__ap_ready;
  wire Mmap2Stream_16__ap_done;
  wire Mmap2Stream_16__ap_idle;
  reg [1:0] Mmap2Stream_16__state;
  wire [63:0] Mmap2Stream_17___n__q0;
  wire [63:0] Mmap2Stream_17___rmem17__q0;
  wire Mmap2Stream_17__ap_start_global__q0;
  wire Mmap2Stream_17__is_done__q0;
  wire Mmap2Stream_17__ap_done_global__q0;
  wire Mmap2Stream_17__ap_start;
  wire Mmap2Stream_17__ap_ready;
  wire Mmap2Stream_17__ap_done;
  wire Mmap2Stream_17__ap_idle;
  reg [1:0] Mmap2Stream_17__state;
  wire [63:0] Mmap2Stream_18___n__q0;
  wire [63:0] Mmap2Stream_18___rmem18__q0;
  wire Mmap2Stream_18__ap_start_global__q0;
  wire Mmap2Stream_18__is_done__q0;
  wire Mmap2Stream_18__ap_done_global__q0;
  wire Mmap2Stream_18__ap_start;
  wire Mmap2Stream_18__ap_ready;
  wire Mmap2Stream_18__ap_done;
  wire Mmap2Stream_18__ap_idle;
  reg [1:0] Mmap2Stream_18__state;
  wire [63:0] Mmap2Stream_19___n__q0;
  wire [63:0] Mmap2Stream_19___rmem19__q0;
  wire Mmap2Stream_19__ap_start_global__q0;
  wire Mmap2Stream_19__is_done__q0;
  wire Mmap2Stream_19__ap_done_global__q0;
  wire Mmap2Stream_19__ap_start;
  wire Mmap2Stream_19__ap_ready;
  wire Mmap2Stream_19__ap_done;
  wire Mmap2Stream_19__ap_idle;
  reg [1:0] Mmap2Stream_19__state;
  wire [63:0] Mmap2Stream_20___n__q0;
  wire [63:0] Mmap2Stream_20___rmem20__q0;
  wire Mmap2Stream_20__ap_start_global__q0;
  wire Mmap2Stream_20__is_done__q0;
  wire Mmap2Stream_20__ap_done_global__q0;
  wire Mmap2Stream_20__ap_start;
  wire Mmap2Stream_20__ap_ready;
  wire Mmap2Stream_20__ap_done;
  wire Mmap2Stream_20__ap_idle;
  reg [1:0] Mmap2Stream_20__state;
  wire [63:0] Mmap2Stream_21___n__q0;
  wire [63:0] Mmap2Stream_21___rmem21__q0;
  wire Mmap2Stream_21__ap_start_global__q0;
  wire Mmap2Stream_21__is_done__q0;
  wire Mmap2Stream_21__ap_done_global__q0;
  wire Mmap2Stream_21__ap_start;
  wire Mmap2Stream_21__ap_ready;
  wire Mmap2Stream_21__ap_done;
  wire Mmap2Stream_21__ap_idle;
  reg [1:0] Mmap2Stream_21__state;
  wire [63:0] Mmap2Stream_22___n__q0;
  wire [63:0] Mmap2Stream_22___rmem22__q0;
  wire Mmap2Stream_22__ap_start_global__q0;
  wire Mmap2Stream_22__is_done__q0;
  wire Mmap2Stream_22__ap_done_global__q0;
  wire Mmap2Stream_22__ap_start;
  wire Mmap2Stream_22__ap_ready;
  wire Mmap2Stream_22__ap_done;
  wire Mmap2Stream_22__ap_idle;
  reg [1:0] Mmap2Stream_22__state;
  wire [63:0] Mmap2Stream_23___n__q0;
  wire [63:0] Mmap2Stream_23___rmem23__q0;
  wire Mmap2Stream_23__ap_start_global__q0;
  wire Mmap2Stream_23__is_done__q0;
  wire Mmap2Stream_23__ap_done_global__q0;
  wire Mmap2Stream_23__ap_start;
  wire Mmap2Stream_23__ap_ready;
  wire Mmap2Stream_23__ap_done;
  wire Mmap2Stream_23__ap_idle;
  reg [1:0] Mmap2Stream_23__state;
  wire [63:0] Mmap2Stream_24___n__q0;
  wire [63:0] Mmap2Stream_24___rmem24__q0;
  wire Mmap2Stream_24__ap_start_global__q0;
  wire Mmap2Stream_24__is_done__q0;
  wire Mmap2Stream_24__ap_done_global__q0;
  wire Mmap2Stream_24__ap_start;
  wire Mmap2Stream_24__ap_ready;
  wire Mmap2Stream_24__ap_done;
  wire Mmap2Stream_24__ap_idle;
  reg [1:0] Mmap2Stream_24__state;
  wire [63:0] Mmap2Stream_25___n__q0;
  wire [63:0] Mmap2Stream_25___rmem25__q0;
  wire Mmap2Stream_25__ap_start_global__q0;
  wire Mmap2Stream_25__is_done__q0;
  wire Mmap2Stream_25__ap_done_global__q0;
  wire Mmap2Stream_25__ap_start;
  wire Mmap2Stream_25__ap_ready;
  wire Mmap2Stream_25__ap_done;
  wire Mmap2Stream_25__ap_idle;
  reg [1:0] Mmap2Stream_25__state;
  wire [63:0] Mmap2Stream_26___n__q0;
  wire [63:0] Mmap2Stream_26___rmem26__q0;
  wire Mmap2Stream_26__ap_start_global__q0;
  wire Mmap2Stream_26__is_done__q0;
  wire Mmap2Stream_26__ap_done_global__q0;
  wire Mmap2Stream_26__ap_start;
  wire Mmap2Stream_26__ap_ready;
  wire Mmap2Stream_26__ap_done;
  wire Mmap2Stream_26__ap_idle;
  reg [1:0] Mmap2Stream_26__state;
  wire [63:0] Mmap2Stream_27___n__q0;
  wire [63:0] Mmap2Stream_27___rmem27__q0;
  wire Mmap2Stream_27__ap_start_global__q0;
  wire Mmap2Stream_27__is_done__q0;
  wire Mmap2Stream_27__ap_done_global__q0;
  wire Mmap2Stream_27__ap_start;
  wire Mmap2Stream_27__ap_ready;
  wire Mmap2Stream_27__ap_done;
  wire Mmap2Stream_27__ap_idle;
  reg [1:0] Mmap2Stream_27__state;
  wire [63:0] Mmap2Stream_28___n__q0;
  wire [63:0] Mmap2Stream_28___rmem28__q0;
  wire Mmap2Stream_28__ap_start_global__q0;
  wire Mmap2Stream_28__is_done__q0;
  wire Mmap2Stream_28__ap_done_global__q0;
  wire Mmap2Stream_28__ap_start;
  wire Mmap2Stream_28__ap_ready;
  wire Mmap2Stream_28__ap_done;
  wire Mmap2Stream_28__ap_idle;
  reg [1:0] Mmap2Stream_28__state;
  wire [63:0] Mmap2Stream_29___n__q0;
  wire [63:0] Mmap2Stream_29___rmem29__q0;
  wire Mmap2Stream_29__ap_start_global__q0;
  wire Mmap2Stream_29__is_done__q0;
  wire Mmap2Stream_29__ap_done_global__q0;
  wire Mmap2Stream_29__ap_start;
  wire Mmap2Stream_29__ap_ready;
  wire Mmap2Stream_29__ap_done;
  wire Mmap2Stream_29__ap_idle;
  reg [1:0] Mmap2Stream_29__state;
  wire [63:0] Stream2Mmap_0___n__q0;
  wire [63:0] Stream2Mmap_0___wmem0__q0;
  wire Stream2Mmap_0__ap_start_global__q0;
  wire Stream2Mmap_0__is_done__q0;
  wire Stream2Mmap_0__ap_done_global__q0;
  wire Stream2Mmap_0__ap_start;
  wire Stream2Mmap_0__ap_ready;
  wire Stream2Mmap_0__ap_done;
  wire Stream2Mmap_0__ap_idle;
  reg [1:0] Stream2Mmap_0__state;
  wire [63:0] yxor_0___n__q0;
  wire yxor_0__ap_start_global__q0;
  wire yxor_0__is_done__q0;
  wire yxor_0__ap_done_global__q0;
  wire yxor_0__ap_start;
  wire yxor_0__ap_ready;
  wire yxor_0__ap_done;
  wire yxor_0__ap_idle;
  reg [1:0] yxor_0__state;
  wire [63:0] yxor_1___n__q0;
  wire yxor_1__ap_start_global__q0;
  wire yxor_1__is_done__q0;
  wire yxor_1__ap_done_global__q0;
  wire yxor_1__ap_start;
  wire yxor_1__ap_ready;
  wire yxor_1__ap_done;
  wire yxor_1__ap_idle;
  reg [1:0] yxor_1__state;
  wire [63:0] yxor_2___n__q0;
  wire yxor_2__ap_start_global__q0;
  wire yxor_2__is_done__q0;
  wire yxor_2__ap_done_global__q0;
  wire yxor_2__ap_start;
  wire yxor_2__ap_ready;
  wire yxor_2__ap_done;
  wire yxor_2__ap_idle;
  reg [1:0] yxor_2__state;
  wire [63:0] yxor_3___n__q0;
  wire yxor_3__ap_start_global__q0;
  wire yxor_3__is_done__q0;
  wire yxor_3__ap_done_global__q0;
  wire yxor_3__ap_start;
  wire yxor_3__ap_ready;
  wire yxor_3__ap_done;
  wire yxor_3__ap_idle;
  reg [1:0] yxor_3__state;
  wire [63:0] yxor_4___n__q0;
  wire yxor_4__ap_start_global__q0;
  wire yxor_4__is_done__q0;
  wire yxor_4__ap_done_global__q0;
  wire yxor_4__ap_start;
  wire yxor_4__ap_ready;
  wire yxor_4__ap_done;
  wire yxor_4__ap_idle;
  reg [1:0] yxor_4__state;
  wire [63:0] yxor_5___n__q0;
  wire yxor_5__ap_start_global__q0;
  wire yxor_5__is_done__q0;
  wire yxor_5__ap_done_global__q0;
  wire yxor_5__ap_start;
  wire yxor_5__ap_ready;
  wire yxor_5__ap_done;
  wire yxor_5__ap_idle;
  reg [1:0] yxor_5__state;
  wire [63:0] yxor_6___n__q0;
  wire yxor_6__ap_start_global__q0;
  wire yxor_6__is_done__q0;
  wire yxor_6__ap_done_global__q0;
  wire yxor_6__ap_start;
  wire yxor_6__ap_ready;
  wire yxor_6__ap_done;
  wire yxor_6__ap_idle;
  reg [1:0] yxor_6__state;
  wire [63:0] yxor_7___n__q0;
  wire yxor_7__ap_start_global__q0;
  wire yxor_7__is_done__q0;
  wire yxor_7__ap_done_global__q0;
  wire yxor_7__ap_start;
  wire yxor_7__ap_ready;
  wire yxor_7__ap_done;
  wire yxor_7__ap_idle;
  reg [1:0] yxor_7__state;
  wire [63:0] yxor_8___n__q0;
  wire yxor_8__ap_start_global__q0;
  wire yxor_8__is_done__q0;
  wire yxor_8__ap_done_global__q0;
  wire yxor_8__ap_start;
  wire yxor_8__ap_ready;
  wire yxor_8__ap_done;
  wire yxor_8__ap_idle;
  reg [1:0] yxor_8__state;
  wire [63:0] yxor_9___n__q0;
  wire yxor_9__ap_start_global__q0;
  wire yxor_9__is_done__q0;
  wire yxor_9__ap_done_global__q0;
  wire yxor_9__ap_start;
  wire yxor_9__ap_ready;
  wire yxor_9__ap_done;
  wire yxor_9__ap_idle;
  reg [1:0] yxor_9__state;
  wire [63:0] yxor_10___n__q0;
  wire yxor_10__ap_start_global__q0;
  wire yxor_10__is_done__q0;
  wire yxor_10__ap_done_global__q0;
  wire yxor_10__ap_start;
  wire yxor_10__ap_ready;
  wire yxor_10__ap_done;
  wire yxor_10__ap_idle;
  reg [1:0] yxor_10__state;
  wire [63:0] yxor_11___n__q0;
  wire yxor_11__ap_start_global__q0;
  wire yxor_11__is_done__q0;
  wire yxor_11__ap_done_global__q0;
  wire yxor_11__ap_start;
  wire yxor_11__ap_ready;
  wire yxor_11__ap_done;
  wire yxor_11__ap_idle;
  reg [1:0] yxor_11__state;
  wire [63:0] yxor_12___n__q0;
  wire yxor_12__ap_start_global__q0;
  wire yxor_12__is_done__q0;
  wire yxor_12__ap_done_global__q0;
  wire yxor_12__ap_start;
  wire yxor_12__ap_ready;
  wire yxor_12__ap_done;
  wire yxor_12__ap_idle;
  reg [1:0] yxor_12__state;
  wire [63:0] yxor_13___n__q0;
  wire yxor_13__ap_start_global__q0;
  wire yxor_13__is_done__q0;
  wire yxor_13__ap_done_global__q0;
  wire yxor_13__ap_start;
  wire yxor_13__ap_ready;
  wire yxor_13__ap_done;
  wire yxor_13__ap_idle;
  reg [1:0] yxor_13__state;
  wire [63:0] yxor_14___n__q0;
  wire yxor_14__ap_start_global__q0;
  wire yxor_14__is_done__q0;
  wire yxor_14__ap_done_global__q0;
  wire yxor_14__ap_start;
  wire yxor_14__ap_ready;
  wire yxor_14__ap_done;
  wire yxor_14__ap_idle;
  reg [1:0] yxor_14__state;
  wire [63:0] yxor_15___n__q0;
  wire yxor_15__ap_start_global__q0;
  wire yxor_15__is_done__q0;
  wire yxor_15__ap_done_global__q0;
  wire yxor_15__ap_start;
  wire yxor_15__ap_ready;
  wire yxor_15__ap_done;
  wire yxor_15__ap_idle;
  reg [1:0] yxor_15__state;
  wire [63:0] yxor_16___n__q0;
  wire yxor_16__ap_start_global__q0;
  wire yxor_16__is_done__q0;
  wire yxor_16__ap_done_global__q0;
  wire yxor_16__ap_start;
  wire yxor_16__ap_ready;
  wire yxor_16__ap_done;
  wire yxor_16__ap_idle;
  reg [1:0] yxor_16__state;
  wire [63:0] yxor_17___n__q0;
  wire yxor_17__ap_start_global__q0;
  wire yxor_17__is_done__q0;
  wire yxor_17__ap_done_global__q0;
  wire yxor_17__ap_start;
  wire yxor_17__ap_ready;
  wire yxor_17__ap_done;
  wire yxor_17__ap_idle;
  reg [1:0] yxor_17__state;
  wire [63:0] yxor_18___n__q0;
  wire yxor_18__ap_start_global__q0;
  wire yxor_18__is_done__q0;
  wire yxor_18__ap_done_global__q0;
  wire yxor_18__ap_start;
  wire yxor_18__ap_ready;
  wire yxor_18__ap_done;
  wire yxor_18__ap_idle;
  reg [1:0] yxor_18__state;
  wire [63:0] yxor_19___n__q0;
  wire yxor_19__ap_start_global__q0;
  wire yxor_19__is_done__q0;
  wire yxor_19__ap_done_global__q0;
  wire yxor_19__ap_start;
  wire yxor_19__ap_ready;
  wire yxor_19__ap_done;
  wire yxor_19__ap_idle;
  reg [1:0] yxor_19__state;
  wire [63:0] yxor_20___n__q0;
  wire yxor_20__ap_start_global__q0;
  wire yxor_20__is_done__q0;
  wire yxor_20__ap_done_global__q0;
  wire yxor_20__ap_start;
  wire yxor_20__ap_ready;
  wire yxor_20__ap_done;
  wire yxor_20__ap_idle;
  reg [1:0] yxor_20__state;
  wire [63:0] yxor_21___n__q0;
  wire yxor_21__ap_start_global__q0;
  wire yxor_21__is_done__q0;
  wire yxor_21__ap_done_global__q0;
  wire yxor_21__ap_start;
  wire yxor_21__ap_ready;
  wire yxor_21__ap_done;
  wire yxor_21__ap_idle;
  reg [1:0] yxor_21__state;
  wire [63:0] yxor_22___n__q0;
  wire yxor_22__ap_start_global__q0;
  wire yxor_22__is_done__q0;
  wire yxor_22__ap_done_global__q0;
  wire yxor_22__ap_start;
  wire yxor_22__ap_ready;
  wire yxor_22__ap_done;
  wire yxor_22__ap_idle;
  reg [1:0] yxor_22__state;
  wire [63:0] yxor_23___n__q0;
  wire yxor_23__ap_start_global__q0;
  wire yxor_23__is_done__q0;
  wire yxor_23__ap_done_global__q0;
  wire yxor_23__ap_start;
  wire yxor_23__ap_ready;
  wire yxor_23__ap_done;
  wire yxor_23__ap_idle;
  reg [1:0] yxor_23__state;
  wire [63:0] yxor_24___n__q0;
  wire yxor_24__ap_start_global__q0;
  wire yxor_24__is_done__q0;
  wire yxor_24__ap_done_global__q0;
  wire yxor_24__ap_start;
  wire yxor_24__ap_ready;
  wire yxor_24__ap_done;
  wire yxor_24__ap_idle;
  reg [1:0] yxor_24__state;
  wire [63:0] yxor_25___n__q0;
  wire yxor_25__ap_start_global__q0;
  wire yxor_25__is_done__q0;
  wire yxor_25__ap_done_global__q0;
  wire yxor_25__ap_start;
  wire yxor_25__ap_ready;
  wire yxor_25__ap_done;
  wire yxor_25__ap_idle;
  reg [1:0] yxor_25__state;
  wire [63:0] yxor_26___n__q0;
  wire yxor_26__ap_start_global__q0;
  wire yxor_26__is_done__q0;
  wire yxor_26__ap_done_global__q0;
  wire yxor_26__ap_start;
  wire yxor_26__ap_ready;
  wire yxor_26__ap_done;
  wire yxor_26__ap_idle;
  reg [1:0] yxor_26__state;
  wire [63:0] yxor_27___n__q0;
  wire yxor_27__ap_start_global__q0;
  wire yxor_27__is_done__q0;
  wire yxor_27__ap_done_global__q0;
  wire yxor_27__ap_start;
  wire yxor_27__ap_ready;
  wire yxor_27__ap_done;
  wire yxor_27__ap_idle;
  reg [1:0] yxor_27__state;
  wire [63:0] yxor_28___n__q0;
  wire yxor_28__ap_start_global__q0;
  wire yxor_28__is_done__q0;
  wire yxor_28__ap_done_global__q0;
  wire yxor_28__ap_start;
  wire yxor_28__ap_ready;
  wire yxor_28__ap_done;
  wire yxor_28__ap_idle;
  reg [1:0] yxor_28__state;
  reg [1:0] tapa_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  wire ap_done__q0;
  assign Mmap2Stream_0___n__q0 = n;
  assign Mmap2Stream_0___rmem0__q0 = rmem0;
  assign Mmap2Stream_0__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_0__is_done__q0 = (Mmap2Stream_0__state == 2'b10);
  assign Mmap2Stream_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_0__state <= 2'b00;
    end else begin
      if(Mmap2Stream_0__state == 2'b00) begin
        if(Mmap2Stream_0__ap_start_global__q0) begin
          Mmap2Stream_0__state <= 2'b01;
        end
      end
      if(Mmap2Stream_0__state == 2'b01) begin
        if(Mmap2Stream_0__ap_ready) begin
          if(Mmap2Stream_0__ap_done) begin
            Mmap2Stream_0__state <= 2'b10;
          end else begin
            Mmap2Stream_0__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_0__state == 2'b11) begin
        if(Mmap2Stream_0__ap_done) begin
          Mmap2Stream_0__state <= 2'b10;
        end
      end
      if(Mmap2Stream_0__state == 2'b10) begin
        if(Mmap2Stream_0__ap_done_global__q0) begin
          Mmap2Stream_0__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_0__ap_start = (Mmap2Stream_0__state == 2'b01);
  assign Mmap2Stream_1___n__q0 = n;
  assign Mmap2Stream_1___rmem1__q0 = rmem1;
  assign Mmap2Stream_1__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_1__is_done__q0 = (Mmap2Stream_1__state == 2'b10);
  assign Mmap2Stream_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_1__state <= 2'b00;
    end else begin
      if(Mmap2Stream_1__state == 2'b00) begin
        if(Mmap2Stream_1__ap_start_global__q0) begin
          Mmap2Stream_1__state <= 2'b01;
        end
      end
      if(Mmap2Stream_1__state == 2'b01) begin
        if(Mmap2Stream_1__ap_ready) begin
          if(Mmap2Stream_1__ap_done) begin
            Mmap2Stream_1__state <= 2'b10;
          end else begin
            Mmap2Stream_1__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_1__state == 2'b11) begin
        if(Mmap2Stream_1__ap_done) begin
          Mmap2Stream_1__state <= 2'b10;
        end
      end
      if(Mmap2Stream_1__state == 2'b10) begin
        if(Mmap2Stream_1__ap_done_global__q0) begin
          Mmap2Stream_1__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_1__ap_start = (Mmap2Stream_1__state == 2'b01);
  assign Mmap2Stream_2___n__q0 = n;
  assign Mmap2Stream_2___rmem2__q0 = rmem2;
  assign Mmap2Stream_2__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_2__is_done__q0 = (Mmap2Stream_2__state == 2'b10);
  assign Mmap2Stream_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_2__state <= 2'b00;
    end else begin
      if(Mmap2Stream_2__state == 2'b00) begin
        if(Mmap2Stream_2__ap_start_global__q0) begin
          Mmap2Stream_2__state <= 2'b01;
        end
      end
      if(Mmap2Stream_2__state == 2'b01) begin
        if(Mmap2Stream_2__ap_ready) begin
          if(Mmap2Stream_2__ap_done) begin
            Mmap2Stream_2__state <= 2'b10;
          end else begin
            Mmap2Stream_2__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_2__state == 2'b11) begin
        if(Mmap2Stream_2__ap_done) begin
          Mmap2Stream_2__state <= 2'b10;
        end
      end
      if(Mmap2Stream_2__state == 2'b10) begin
        if(Mmap2Stream_2__ap_done_global__q0) begin
          Mmap2Stream_2__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_2__ap_start = (Mmap2Stream_2__state == 2'b01);
  assign Mmap2Stream_3___n__q0 = n;
  assign Mmap2Stream_3___rmem3__q0 = rmem3;
  assign Mmap2Stream_3__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_3__is_done__q0 = (Mmap2Stream_3__state == 2'b10);
  assign Mmap2Stream_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_3__state <= 2'b00;
    end else begin
      if(Mmap2Stream_3__state == 2'b00) begin
        if(Mmap2Stream_3__ap_start_global__q0) begin
          Mmap2Stream_3__state <= 2'b01;
        end
      end
      if(Mmap2Stream_3__state == 2'b01) begin
        if(Mmap2Stream_3__ap_ready) begin
          if(Mmap2Stream_3__ap_done) begin
            Mmap2Stream_3__state <= 2'b10;
          end else begin
            Mmap2Stream_3__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_3__state == 2'b11) begin
        if(Mmap2Stream_3__ap_done) begin
          Mmap2Stream_3__state <= 2'b10;
        end
      end
      if(Mmap2Stream_3__state == 2'b10) begin
        if(Mmap2Stream_3__ap_done_global__q0) begin
          Mmap2Stream_3__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_3__ap_start = (Mmap2Stream_3__state == 2'b01);
  assign Mmap2Stream_4___n__q0 = n;
  assign Mmap2Stream_4___rmem4__q0 = rmem4;
  assign Mmap2Stream_4__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_4__is_done__q0 = (Mmap2Stream_4__state == 2'b10);
  assign Mmap2Stream_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_4__state <= 2'b00;
    end else begin
      if(Mmap2Stream_4__state == 2'b00) begin
        if(Mmap2Stream_4__ap_start_global__q0) begin
          Mmap2Stream_4__state <= 2'b01;
        end
      end
      if(Mmap2Stream_4__state == 2'b01) begin
        if(Mmap2Stream_4__ap_ready) begin
          if(Mmap2Stream_4__ap_done) begin
            Mmap2Stream_4__state <= 2'b10;
          end else begin
            Mmap2Stream_4__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_4__state == 2'b11) begin
        if(Mmap2Stream_4__ap_done) begin
          Mmap2Stream_4__state <= 2'b10;
        end
      end
      if(Mmap2Stream_4__state == 2'b10) begin
        if(Mmap2Stream_4__ap_done_global__q0) begin
          Mmap2Stream_4__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_4__ap_start = (Mmap2Stream_4__state == 2'b01);
  assign Mmap2Stream_5___n__q0 = n;
  assign Mmap2Stream_5___rmem5__q0 = rmem5;
  assign Mmap2Stream_5__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_5__is_done__q0 = (Mmap2Stream_5__state == 2'b10);
  assign Mmap2Stream_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_5__state <= 2'b00;
    end else begin
      if(Mmap2Stream_5__state == 2'b00) begin
        if(Mmap2Stream_5__ap_start_global__q0) begin
          Mmap2Stream_5__state <= 2'b01;
        end
      end
      if(Mmap2Stream_5__state == 2'b01) begin
        if(Mmap2Stream_5__ap_ready) begin
          if(Mmap2Stream_5__ap_done) begin
            Mmap2Stream_5__state <= 2'b10;
          end else begin
            Mmap2Stream_5__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_5__state == 2'b11) begin
        if(Mmap2Stream_5__ap_done) begin
          Mmap2Stream_5__state <= 2'b10;
        end
      end
      if(Mmap2Stream_5__state == 2'b10) begin
        if(Mmap2Stream_5__ap_done_global__q0) begin
          Mmap2Stream_5__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_5__ap_start = (Mmap2Stream_5__state == 2'b01);
  assign Mmap2Stream_6___n__q0 = n;
  assign Mmap2Stream_6___rmem6__q0 = rmem6;
  assign Mmap2Stream_6__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_6__is_done__q0 = (Mmap2Stream_6__state == 2'b10);
  assign Mmap2Stream_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_6__state <= 2'b00;
    end else begin
      if(Mmap2Stream_6__state == 2'b00) begin
        if(Mmap2Stream_6__ap_start_global__q0) begin
          Mmap2Stream_6__state <= 2'b01;
        end
      end
      if(Mmap2Stream_6__state == 2'b01) begin
        if(Mmap2Stream_6__ap_ready) begin
          if(Mmap2Stream_6__ap_done) begin
            Mmap2Stream_6__state <= 2'b10;
          end else begin
            Mmap2Stream_6__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_6__state == 2'b11) begin
        if(Mmap2Stream_6__ap_done) begin
          Mmap2Stream_6__state <= 2'b10;
        end
      end
      if(Mmap2Stream_6__state == 2'b10) begin
        if(Mmap2Stream_6__ap_done_global__q0) begin
          Mmap2Stream_6__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_6__ap_start = (Mmap2Stream_6__state == 2'b01);
  assign Mmap2Stream_7___n__q0 = n;
  assign Mmap2Stream_7___rmem7__q0 = rmem7;
  assign Mmap2Stream_7__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_7__is_done__q0 = (Mmap2Stream_7__state == 2'b10);
  assign Mmap2Stream_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_7__state <= 2'b00;
    end else begin
      if(Mmap2Stream_7__state == 2'b00) begin
        if(Mmap2Stream_7__ap_start_global__q0) begin
          Mmap2Stream_7__state <= 2'b01;
        end
      end
      if(Mmap2Stream_7__state == 2'b01) begin
        if(Mmap2Stream_7__ap_ready) begin
          if(Mmap2Stream_7__ap_done) begin
            Mmap2Stream_7__state <= 2'b10;
          end else begin
            Mmap2Stream_7__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_7__state == 2'b11) begin
        if(Mmap2Stream_7__ap_done) begin
          Mmap2Stream_7__state <= 2'b10;
        end
      end
      if(Mmap2Stream_7__state == 2'b10) begin
        if(Mmap2Stream_7__ap_done_global__q0) begin
          Mmap2Stream_7__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_7__ap_start = (Mmap2Stream_7__state == 2'b01);
  assign Mmap2Stream_8___n__q0 = n;
  assign Mmap2Stream_8___rmem8__q0 = rmem8;
  assign Mmap2Stream_8__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_8__is_done__q0 = (Mmap2Stream_8__state == 2'b10);
  assign Mmap2Stream_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_8__state <= 2'b00;
    end else begin
      if(Mmap2Stream_8__state == 2'b00) begin
        if(Mmap2Stream_8__ap_start_global__q0) begin
          Mmap2Stream_8__state <= 2'b01;
        end
      end
      if(Mmap2Stream_8__state == 2'b01) begin
        if(Mmap2Stream_8__ap_ready) begin
          if(Mmap2Stream_8__ap_done) begin
            Mmap2Stream_8__state <= 2'b10;
          end else begin
            Mmap2Stream_8__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_8__state == 2'b11) begin
        if(Mmap2Stream_8__ap_done) begin
          Mmap2Stream_8__state <= 2'b10;
        end
      end
      if(Mmap2Stream_8__state == 2'b10) begin
        if(Mmap2Stream_8__ap_done_global__q0) begin
          Mmap2Stream_8__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_8__ap_start = (Mmap2Stream_8__state == 2'b01);
  assign Mmap2Stream_9___n__q0 = n;
  assign Mmap2Stream_9___rmem9__q0 = rmem9;
  assign Mmap2Stream_9__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_9__is_done__q0 = (Mmap2Stream_9__state == 2'b10);
  assign Mmap2Stream_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_9__state <= 2'b00;
    end else begin
      if(Mmap2Stream_9__state == 2'b00) begin
        if(Mmap2Stream_9__ap_start_global__q0) begin
          Mmap2Stream_9__state <= 2'b01;
        end
      end
      if(Mmap2Stream_9__state == 2'b01) begin
        if(Mmap2Stream_9__ap_ready) begin
          if(Mmap2Stream_9__ap_done) begin
            Mmap2Stream_9__state <= 2'b10;
          end else begin
            Mmap2Stream_9__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_9__state == 2'b11) begin
        if(Mmap2Stream_9__ap_done) begin
          Mmap2Stream_9__state <= 2'b10;
        end
      end
      if(Mmap2Stream_9__state == 2'b10) begin
        if(Mmap2Stream_9__ap_done_global__q0) begin
          Mmap2Stream_9__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_9__ap_start = (Mmap2Stream_9__state == 2'b01);
  assign Mmap2Stream_10___n__q0 = n;
  assign Mmap2Stream_10___rmem10__q0 = rmem10;
  assign Mmap2Stream_10__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_10__is_done__q0 = (Mmap2Stream_10__state == 2'b10);
  assign Mmap2Stream_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_10__state <= 2'b00;
    end else begin
      if(Mmap2Stream_10__state == 2'b00) begin
        if(Mmap2Stream_10__ap_start_global__q0) begin
          Mmap2Stream_10__state <= 2'b01;
        end
      end
      if(Mmap2Stream_10__state == 2'b01) begin
        if(Mmap2Stream_10__ap_ready) begin
          if(Mmap2Stream_10__ap_done) begin
            Mmap2Stream_10__state <= 2'b10;
          end else begin
            Mmap2Stream_10__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_10__state == 2'b11) begin
        if(Mmap2Stream_10__ap_done) begin
          Mmap2Stream_10__state <= 2'b10;
        end
      end
      if(Mmap2Stream_10__state == 2'b10) begin
        if(Mmap2Stream_10__ap_done_global__q0) begin
          Mmap2Stream_10__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_10__ap_start = (Mmap2Stream_10__state == 2'b01);
  assign Mmap2Stream_11___n__q0 = n;
  assign Mmap2Stream_11___rmem11__q0 = rmem11;
  assign Mmap2Stream_11__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_11__is_done__q0 = (Mmap2Stream_11__state == 2'b10);
  assign Mmap2Stream_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_11__state <= 2'b00;
    end else begin
      if(Mmap2Stream_11__state == 2'b00) begin
        if(Mmap2Stream_11__ap_start_global__q0) begin
          Mmap2Stream_11__state <= 2'b01;
        end
      end
      if(Mmap2Stream_11__state == 2'b01) begin
        if(Mmap2Stream_11__ap_ready) begin
          if(Mmap2Stream_11__ap_done) begin
            Mmap2Stream_11__state <= 2'b10;
          end else begin
            Mmap2Stream_11__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_11__state == 2'b11) begin
        if(Mmap2Stream_11__ap_done) begin
          Mmap2Stream_11__state <= 2'b10;
        end
      end
      if(Mmap2Stream_11__state == 2'b10) begin
        if(Mmap2Stream_11__ap_done_global__q0) begin
          Mmap2Stream_11__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_11__ap_start = (Mmap2Stream_11__state == 2'b01);
  assign Mmap2Stream_12___n__q0 = n;
  assign Mmap2Stream_12___rmem12__q0 = rmem12;
  assign Mmap2Stream_12__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_12__is_done__q0 = (Mmap2Stream_12__state == 2'b10);
  assign Mmap2Stream_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_12__state <= 2'b00;
    end else begin
      if(Mmap2Stream_12__state == 2'b00) begin
        if(Mmap2Stream_12__ap_start_global__q0) begin
          Mmap2Stream_12__state <= 2'b01;
        end
      end
      if(Mmap2Stream_12__state == 2'b01) begin
        if(Mmap2Stream_12__ap_ready) begin
          if(Mmap2Stream_12__ap_done) begin
            Mmap2Stream_12__state <= 2'b10;
          end else begin
            Mmap2Stream_12__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_12__state == 2'b11) begin
        if(Mmap2Stream_12__ap_done) begin
          Mmap2Stream_12__state <= 2'b10;
        end
      end
      if(Mmap2Stream_12__state == 2'b10) begin
        if(Mmap2Stream_12__ap_done_global__q0) begin
          Mmap2Stream_12__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_12__ap_start = (Mmap2Stream_12__state == 2'b01);
  assign Mmap2Stream_13___n__q0 = n;
  assign Mmap2Stream_13___rmem13__q0 = rmem13;
  assign Mmap2Stream_13__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_13__is_done__q0 = (Mmap2Stream_13__state == 2'b10);
  assign Mmap2Stream_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_13__state <= 2'b00;
    end else begin
      if(Mmap2Stream_13__state == 2'b00) begin
        if(Mmap2Stream_13__ap_start_global__q0) begin
          Mmap2Stream_13__state <= 2'b01;
        end
      end
      if(Mmap2Stream_13__state == 2'b01) begin
        if(Mmap2Stream_13__ap_ready) begin
          if(Mmap2Stream_13__ap_done) begin
            Mmap2Stream_13__state <= 2'b10;
          end else begin
            Mmap2Stream_13__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_13__state == 2'b11) begin
        if(Mmap2Stream_13__ap_done) begin
          Mmap2Stream_13__state <= 2'b10;
        end
      end
      if(Mmap2Stream_13__state == 2'b10) begin
        if(Mmap2Stream_13__ap_done_global__q0) begin
          Mmap2Stream_13__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_13__ap_start = (Mmap2Stream_13__state == 2'b01);
  assign Mmap2Stream_14___n__q0 = n;
  assign Mmap2Stream_14___rmem14__q0 = rmem14;
  assign Mmap2Stream_14__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_14__is_done__q0 = (Mmap2Stream_14__state == 2'b10);
  assign Mmap2Stream_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_14__state <= 2'b00;
    end else begin
      if(Mmap2Stream_14__state == 2'b00) begin
        if(Mmap2Stream_14__ap_start_global__q0) begin
          Mmap2Stream_14__state <= 2'b01;
        end
      end
      if(Mmap2Stream_14__state == 2'b01) begin
        if(Mmap2Stream_14__ap_ready) begin
          if(Mmap2Stream_14__ap_done) begin
            Mmap2Stream_14__state <= 2'b10;
          end else begin
            Mmap2Stream_14__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_14__state == 2'b11) begin
        if(Mmap2Stream_14__ap_done) begin
          Mmap2Stream_14__state <= 2'b10;
        end
      end
      if(Mmap2Stream_14__state == 2'b10) begin
        if(Mmap2Stream_14__ap_done_global__q0) begin
          Mmap2Stream_14__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_14__ap_start = (Mmap2Stream_14__state == 2'b01);
  assign Mmap2Stream_15___n__q0 = n;
  assign Mmap2Stream_15___rmem15__q0 = rmem15;
  assign Mmap2Stream_15__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_15__is_done__q0 = (Mmap2Stream_15__state == 2'b10);
  assign Mmap2Stream_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_15__state <= 2'b00;
    end else begin
      if(Mmap2Stream_15__state == 2'b00) begin
        if(Mmap2Stream_15__ap_start_global__q0) begin
          Mmap2Stream_15__state <= 2'b01;
        end
      end
      if(Mmap2Stream_15__state == 2'b01) begin
        if(Mmap2Stream_15__ap_ready) begin
          if(Mmap2Stream_15__ap_done) begin
            Mmap2Stream_15__state <= 2'b10;
          end else begin
            Mmap2Stream_15__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_15__state == 2'b11) begin
        if(Mmap2Stream_15__ap_done) begin
          Mmap2Stream_15__state <= 2'b10;
        end
      end
      if(Mmap2Stream_15__state == 2'b10) begin
        if(Mmap2Stream_15__ap_done_global__q0) begin
          Mmap2Stream_15__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_15__ap_start = (Mmap2Stream_15__state == 2'b01);
  assign Mmap2Stream_16___n__q0 = n;
  assign Mmap2Stream_16___rmem16__q0 = rmem16;
  assign Mmap2Stream_16__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_16__is_done__q0 = (Mmap2Stream_16__state == 2'b10);
  assign Mmap2Stream_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_16__state <= 2'b00;
    end else begin
      if(Mmap2Stream_16__state == 2'b00) begin
        if(Mmap2Stream_16__ap_start_global__q0) begin
          Mmap2Stream_16__state <= 2'b01;
        end
      end
      if(Mmap2Stream_16__state == 2'b01) begin
        if(Mmap2Stream_16__ap_ready) begin
          if(Mmap2Stream_16__ap_done) begin
            Mmap2Stream_16__state <= 2'b10;
          end else begin
            Mmap2Stream_16__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_16__state == 2'b11) begin
        if(Mmap2Stream_16__ap_done) begin
          Mmap2Stream_16__state <= 2'b10;
        end
      end
      if(Mmap2Stream_16__state == 2'b10) begin
        if(Mmap2Stream_16__ap_done_global__q0) begin
          Mmap2Stream_16__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_16__ap_start = (Mmap2Stream_16__state == 2'b01);
  assign Mmap2Stream_17___n__q0 = n;
  assign Mmap2Stream_17___rmem17__q0 = rmem17;
  assign Mmap2Stream_17__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_17__is_done__q0 = (Mmap2Stream_17__state == 2'b10);
  assign Mmap2Stream_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_17__state <= 2'b00;
    end else begin
      if(Mmap2Stream_17__state == 2'b00) begin
        if(Mmap2Stream_17__ap_start_global__q0) begin
          Mmap2Stream_17__state <= 2'b01;
        end
      end
      if(Mmap2Stream_17__state == 2'b01) begin
        if(Mmap2Stream_17__ap_ready) begin
          if(Mmap2Stream_17__ap_done) begin
            Mmap2Stream_17__state <= 2'b10;
          end else begin
            Mmap2Stream_17__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_17__state == 2'b11) begin
        if(Mmap2Stream_17__ap_done) begin
          Mmap2Stream_17__state <= 2'b10;
        end
      end
      if(Mmap2Stream_17__state == 2'b10) begin
        if(Mmap2Stream_17__ap_done_global__q0) begin
          Mmap2Stream_17__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_17__ap_start = (Mmap2Stream_17__state == 2'b01);
  assign Mmap2Stream_18___n__q0 = n;
  assign Mmap2Stream_18___rmem18__q0 = rmem18;
  assign Mmap2Stream_18__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_18__is_done__q0 = (Mmap2Stream_18__state == 2'b10);
  assign Mmap2Stream_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_18__state <= 2'b00;
    end else begin
      if(Mmap2Stream_18__state == 2'b00) begin
        if(Mmap2Stream_18__ap_start_global__q0) begin
          Mmap2Stream_18__state <= 2'b01;
        end
      end
      if(Mmap2Stream_18__state == 2'b01) begin
        if(Mmap2Stream_18__ap_ready) begin
          if(Mmap2Stream_18__ap_done) begin
            Mmap2Stream_18__state <= 2'b10;
          end else begin
            Mmap2Stream_18__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_18__state == 2'b11) begin
        if(Mmap2Stream_18__ap_done) begin
          Mmap2Stream_18__state <= 2'b10;
        end
      end
      if(Mmap2Stream_18__state == 2'b10) begin
        if(Mmap2Stream_18__ap_done_global__q0) begin
          Mmap2Stream_18__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_18__ap_start = (Mmap2Stream_18__state == 2'b01);
  assign Mmap2Stream_19___n__q0 = n;
  assign Mmap2Stream_19___rmem19__q0 = rmem19;
  assign Mmap2Stream_19__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_19__is_done__q0 = (Mmap2Stream_19__state == 2'b10);
  assign Mmap2Stream_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_19__state <= 2'b00;
    end else begin
      if(Mmap2Stream_19__state == 2'b00) begin
        if(Mmap2Stream_19__ap_start_global__q0) begin
          Mmap2Stream_19__state <= 2'b01;
        end
      end
      if(Mmap2Stream_19__state == 2'b01) begin
        if(Mmap2Stream_19__ap_ready) begin
          if(Mmap2Stream_19__ap_done) begin
            Mmap2Stream_19__state <= 2'b10;
          end else begin
            Mmap2Stream_19__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_19__state == 2'b11) begin
        if(Mmap2Stream_19__ap_done) begin
          Mmap2Stream_19__state <= 2'b10;
        end
      end
      if(Mmap2Stream_19__state == 2'b10) begin
        if(Mmap2Stream_19__ap_done_global__q0) begin
          Mmap2Stream_19__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_19__ap_start = (Mmap2Stream_19__state == 2'b01);
  assign Mmap2Stream_20___n__q0 = n;
  assign Mmap2Stream_20___rmem20__q0 = rmem20;
  assign Mmap2Stream_20__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_20__is_done__q0 = (Mmap2Stream_20__state == 2'b10);
  assign Mmap2Stream_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_20__state <= 2'b00;
    end else begin
      if(Mmap2Stream_20__state == 2'b00) begin
        if(Mmap2Stream_20__ap_start_global__q0) begin
          Mmap2Stream_20__state <= 2'b01;
        end
      end
      if(Mmap2Stream_20__state == 2'b01) begin
        if(Mmap2Stream_20__ap_ready) begin
          if(Mmap2Stream_20__ap_done) begin
            Mmap2Stream_20__state <= 2'b10;
          end else begin
            Mmap2Stream_20__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_20__state == 2'b11) begin
        if(Mmap2Stream_20__ap_done) begin
          Mmap2Stream_20__state <= 2'b10;
        end
      end
      if(Mmap2Stream_20__state == 2'b10) begin
        if(Mmap2Stream_20__ap_done_global__q0) begin
          Mmap2Stream_20__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_20__ap_start = (Mmap2Stream_20__state == 2'b01);
  assign Mmap2Stream_21___n__q0 = n;
  assign Mmap2Stream_21___rmem21__q0 = rmem21;
  assign Mmap2Stream_21__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_21__is_done__q0 = (Mmap2Stream_21__state == 2'b10);
  assign Mmap2Stream_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_21__state <= 2'b00;
    end else begin
      if(Mmap2Stream_21__state == 2'b00) begin
        if(Mmap2Stream_21__ap_start_global__q0) begin
          Mmap2Stream_21__state <= 2'b01;
        end
      end
      if(Mmap2Stream_21__state == 2'b01) begin
        if(Mmap2Stream_21__ap_ready) begin
          if(Mmap2Stream_21__ap_done) begin
            Mmap2Stream_21__state <= 2'b10;
          end else begin
            Mmap2Stream_21__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_21__state == 2'b11) begin
        if(Mmap2Stream_21__ap_done) begin
          Mmap2Stream_21__state <= 2'b10;
        end
      end
      if(Mmap2Stream_21__state == 2'b10) begin
        if(Mmap2Stream_21__ap_done_global__q0) begin
          Mmap2Stream_21__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_21__ap_start = (Mmap2Stream_21__state == 2'b01);
  assign Mmap2Stream_22___n__q0 = n;
  assign Mmap2Stream_22___rmem22__q0 = rmem22;
  assign Mmap2Stream_22__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_22__is_done__q0 = (Mmap2Stream_22__state == 2'b10);
  assign Mmap2Stream_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_22__state <= 2'b00;
    end else begin
      if(Mmap2Stream_22__state == 2'b00) begin
        if(Mmap2Stream_22__ap_start_global__q0) begin
          Mmap2Stream_22__state <= 2'b01;
        end
      end
      if(Mmap2Stream_22__state == 2'b01) begin
        if(Mmap2Stream_22__ap_ready) begin
          if(Mmap2Stream_22__ap_done) begin
            Mmap2Stream_22__state <= 2'b10;
          end else begin
            Mmap2Stream_22__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_22__state == 2'b11) begin
        if(Mmap2Stream_22__ap_done) begin
          Mmap2Stream_22__state <= 2'b10;
        end
      end
      if(Mmap2Stream_22__state == 2'b10) begin
        if(Mmap2Stream_22__ap_done_global__q0) begin
          Mmap2Stream_22__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_22__ap_start = (Mmap2Stream_22__state == 2'b01);
  assign Mmap2Stream_23___n__q0 = n;
  assign Mmap2Stream_23___rmem23__q0 = rmem23;
  assign Mmap2Stream_23__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_23__is_done__q0 = (Mmap2Stream_23__state == 2'b10);
  assign Mmap2Stream_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_23__state <= 2'b00;
    end else begin
      if(Mmap2Stream_23__state == 2'b00) begin
        if(Mmap2Stream_23__ap_start_global__q0) begin
          Mmap2Stream_23__state <= 2'b01;
        end
      end
      if(Mmap2Stream_23__state == 2'b01) begin
        if(Mmap2Stream_23__ap_ready) begin
          if(Mmap2Stream_23__ap_done) begin
            Mmap2Stream_23__state <= 2'b10;
          end else begin
            Mmap2Stream_23__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_23__state == 2'b11) begin
        if(Mmap2Stream_23__ap_done) begin
          Mmap2Stream_23__state <= 2'b10;
        end
      end
      if(Mmap2Stream_23__state == 2'b10) begin
        if(Mmap2Stream_23__ap_done_global__q0) begin
          Mmap2Stream_23__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_23__ap_start = (Mmap2Stream_23__state == 2'b01);
  assign Mmap2Stream_24___n__q0 = n;
  assign Mmap2Stream_24___rmem24__q0 = rmem24;
  assign Mmap2Stream_24__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_24__is_done__q0 = (Mmap2Stream_24__state == 2'b10);
  assign Mmap2Stream_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_24__state <= 2'b00;
    end else begin
      if(Mmap2Stream_24__state == 2'b00) begin
        if(Mmap2Stream_24__ap_start_global__q0) begin
          Mmap2Stream_24__state <= 2'b01;
        end
      end
      if(Mmap2Stream_24__state == 2'b01) begin
        if(Mmap2Stream_24__ap_ready) begin
          if(Mmap2Stream_24__ap_done) begin
            Mmap2Stream_24__state <= 2'b10;
          end else begin
            Mmap2Stream_24__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_24__state == 2'b11) begin
        if(Mmap2Stream_24__ap_done) begin
          Mmap2Stream_24__state <= 2'b10;
        end
      end
      if(Mmap2Stream_24__state == 2'b10) begin
        if(Mmap2Stream_24__ap_done_global__q0) begin
          Mmap2Stream_24__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_24__ap_start = (Mmap2Stream_24__state == 2'b01);
  assign Mmap2Stream_25___n__q0 = n;
  assign Mmap2Stream_25___rmem25__q0 = rmem25;
  assign Mmap2Stream_25__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_25__is_done__q0 = (Mmap2Stream_25__state == 2'b10);
  assign Mmap2Stream_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_25__state <= 2'b00;
    end else begin
      if(Mmap2Stream_25__state == 2'b00) begin
        if(Mmap2Stream_25__ap_start_global__q0) begin
          Mmap2Stream_25__state <= 2'b01;
        end
      end
      if(Mmap2Stream_25__state == 2'b01) begin
        if(Mmap2Stream_25__ap_ready) begin
          if(Mmap2Stream_25__ap_done) begin
            Mmap2Stream_25__state <= 2'b10;
          end else begin
            Mmap2Stream_25__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_25__state == 2'b11) begin
        if(Mmap2Stream_25__ap_done) begin
          Mmap2Stream_25__state <= 2'b10;
        end
      end
      if(Mmap2Stream_25__state == 2'b10) begin
        if(Mmap2Stream_25__ap_done_global__q0) begin
          Mmap2Stream_25__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_25__ap_start = (Mmap2Stream_25__state == 2'b01);
  assign Mmap2Stream_26___n__q0 = n;
  assign Mmap2Stream_26___rmem26__q0 = rmem26;
  assign Mmap2Stream_26__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_26__is_done__q0 = (Mmap2Stream_26__state == 2'b10);
  assign Mmap2Stream_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_26__state <= 2'b00;
    end else begin
      if(Mmap2Stream_26__state == 2'b00) begin
        if(Mmap2Stream_26__ap_start_global__q0) begin
          Mmap2Stream_26__state <= 2'b01;
        end
      end
      if(Mmap2Stream_26__state == 2'b01) begin
        if(Mmap2Stream_26__ap_ready) begin
          if(Mmap2Stream_26__ap_done) begin
            Mmap2Stream_26__state <= 2'b10;
          end else begin
            Mmap2Stream_26__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_26__state == 2'b11) begin
        if(Mmap2Stream_26__ap_done) begin
          Mmap2Stream_26__state <= 2'b10;
        end
      end
      if(Mmap2Stream_26__state == 2'b10) begin
        if(Mmap2Stream_26__ap_done_global__q0) begin
          Mmap2Stream_26__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_26__ap_start = (Mmap2Stream_26__state == 2'b01);
  assign Mmap2Stream_27___n__q0 = n;
  assign Mmap2Stream_27___rmem27__q0 = rmem27;
  assign Mmap2Stream_27__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_27__is_done__q0 = (Mmap2Stream_27__state == 2'b10);
  assign Mmap2Stream_27__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_27__state <= 2'b00;
    end else begin
      if(Mmap2Stream_27__state == 2'b00) begin
        if(Mmap2Stream_27__ap_start_global__q0) begin
          Mmap2Stream_27__state <= 2'b01;
        end
      end
      if(Mmap2Stream_27__state == 2'b01) begin
        if(Mmap2Stream_27__ap_ready) begin
          if(Mmap2Stream_27__ap_done) begin
            Mmap2Stream_27__state <= 2'b10;
          end else begin
            Mmap2Stream_27__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_27__state == 2'b11) begin
        if(Mmap2Stream_27__ap_done) begin
          Mmap2Stream_27__state <= 2'b10;
        end
      end
      if(Mmap2Stream_27__state == 2'b10) begin
        if(Mmap2Stream_27__ap_done_global__q0) begin
          Mmap2Stream_27__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_27__ap_start = (Mmap2Stream_27__state == 2'b01);
  assign Mmap2Stream_28___n__q0 = n;
  assign Mmap2Stream_28___rmem28__q0 = rmem28;
  assign Mmap2Stream_28__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_28__is_done__q0 = (Mmap2Stream_28__state == 2'b10);
  assign Mmap2Stream_28__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_28__state <= 2'b00;
    end else begin
      if(Mmap2Stream_28__state == 2'b00) begin
        if(Mmap2Stream_28__ap_start_global__q0) begin
          Mmap2Stream_28__state <= 2'b01;
        end
      end
      if(Mmap2Stream_28__state == 2'b01) begin
        if(Mmap2Stream_28__ap_ready) begin
          if(Mmap2Stream_28__ap_done) begin
            Mmap2Stream_28__state <= 2'b10;
          end else begin
            Mmap2Stream_28__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_28__state == 2'b11) begin
        if(Mmap2Stream_28__ap_done) begin
          Mmap2Stream_28__state <= 2'b10;
        end
      end
      if(Mmap2Stream_28__state == 2'b10) begin
        if(Mmap2Stream_28__ap_done_global__q0) begin
          Mmap2Stream_28__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_28__ap_start = (Mmap2Stream_28__state == 2'b01);
  assign Mmap2Stream_29___n__q0 = n;
  assign Mmap2Stream_29___rmem29__q0 = rmem29;
  assign Mmap2Stream_29__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_29__is_done__q0 = (Mmap2Stream_29__state == 2'b10);
  assign Mmap2Stream_29__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_29__state <= 2'b00;
    end else begin
      if(Mmap2Stream_29__state == 2'b00) begin
        if(Mmap2Stream_29__ap_start_global__q0) begin
          Mmap2Stream_29__state <= 2'b01;
        end
      end
      if(Mmap2Stream_29__state == 2'b01) begin
        if(Mmap2Stream_29__ap_ready) begin
          if(Mmap2Stream_29__ap_done) begin
            Mmap2Stream_29__state <= 2'b10;
          end else begin
            Mmap2Stream_29__state <= 2'b11;
          end
        end
      end
      if(Mmap2Stream_29__state == 2'b11) begin
        if(Mmap2Stream_29__ap_done) begin
          Mmap2Stream_29__state <= 2'b10;
        end
      end
      if(Mmap2Stream_29__state == 2'b10) begin
        if(Mmap2Stream_29__ap_done_global__q0) begin
          Mmap2Stream_29__state <= 2'b00;
        end
      end
    end
  end

  assign Mmap2Stream_29__ap_start = (Mmap2Stream_29__state == 2'b01);
  assign Stream2Mmap_0___n__q0 = n;
  assign Stream2Mmap_0___wmem0__q0 = wmem0;
  assign Stream2Mmap_0__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_0__is_done__q0 = (Stream2Mmap_0__state == 2'b10);
  assign Stream2Mmap_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_0__state <= 2'b00;
    end else begin
      if(Stream2Mmap_0__state == 2'b00) begin
        if(Stream2Mmap_0__ap_start_global__q0) begin
          Stream2Mmap_0__state <= 2'b01;
        end
      end
      if(Stream2Mmap_0__state == 2'b01) begin
        if(Stream2Mmap_0__ap_ready) begin
          if(Stream2Mmap_0__ap_done) begin
            Stream2Mmap_0__state <= 2'b10;
          end else begin
            Stream2Mmap_0__state <= 2'b11;
          end
        end
      end
      if(Stream2Mmap_0__state == 2'b11) begin
        if(Stream2Mmap_0__ap_done) begin
          Stream2Mmap_0__state <= 2'b10;
        end
      end
      if(Stream2Mmap_0__state == 2'b10) begin
        if(Stream2Mmap_0__ap_done_global__q0) begin
          Stream2Mmap_0__state <= 2'b00;
        end
      end
    end
  end

  assign Stream2Mmap_0__ap_start = (Stream2Mmap_0__state == 2'b01);
  assign yxor_0___n__q0 = n;
  assign yxor_0__ap_start_global__q0 = ap_start__q0;
  assign yxor_0__is_done__q0 = (yxor_0__state == 2'b10);
  assign yxor_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_0__state <= 2'b00;
    end else begin
      if(yxor_0__state == 2'b00) begin
        if(yxor_0__ap_start_global__q0) begin
          yxor_0__state <= 2'b01;
        end
      end
      if(yxor_0__state == 2'b01) begin
        if(yxor_0__ap_ready) begin
          if(yxor_0__ap_done) begin
            yxor_0__state <= 2'b10;
          end else begin
            yxor_0__state <= 2'b11;
          end
        end
      end
      if(yxor_0__state == 2'b11) begin
        if(yxor_0__ap_done) begin
          yxor_0__state <= 2'b10;
        end
      end
      if(yxor_0__state == 2'b10) begin
        if(yxor_0__ap_done_global__q0) begin
          yxor_0__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_0__ap_start = (yxor_0__state == 2'b01);
  assign yxor_1___n__q0 = n;
  assign yxor_1__ap_start_global__q0 = ap_start__q0;
  assign yxor_1__is_done__q0 = (yxor_1__state == 2'b10);
  assign yxor_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_1__state <= 2'b00;
    end else begin
      if(yxor_1__state == 2'b00) begin
        if(yxor_1__ap_start_global__q0) begin
          yxor_1__state <= 2'b01;
        end
      end
      if(yxor_1__state == 2'b01) begin
        if(yxor_1__ap_ready) begin
          if(yxor_1__ap_done) begin
            yxor_1__state <= 2'b10;
          end else begin
            yxor_1__state <= 2'b11;
          end
        end
      end
      if(yxor_1__state == 2'b11) begin
        if(yxor_1__ap_done) begin
          yxor_1__state <= 2'b10;
        end
      end
      if(yxor_1__state == 2'b10) begin
        if(yxor_1__ap_done_global__q0) begin
          yxor_1__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_1__ap_start = (yxor_1__state == 2'b01);
  assign yxor_2___n__q0 = n;
  assign yxor_2__ap_start_global__q0 = ap_start__q0;
  assign yxor_2__is_done__q0 = (yxor_2__state == 2'b10);
  assign yxor_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_2__state <= 2'b00;
    end else begin
      if(yxor_2__state == 2'b00) begin
        if(yxor_2__ap_start_global__q0) begin
          yxor_2__state <= 2'b01;
        end
      end
      if(yxor_2__state == 2'b01) begin
        if(yxor_2__ap_ready) begin
          if(yxor_2__ap_done) begin
            yxor_2__state <= 2'b10;
          end else begin
            yxor_2__state <= 2'b11;
          end
        end
      end
      if(yxor_2__state == 2'b11) begin
        if(yxor_2__ap_done) begin
          yxor_2__state <= 2'b10;
        end
      end
      if(yxor_2__state == 2'b10) begin
        if(yxor_2__ap_done_global__q0) begin
          yxor_2__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_2__ap_start = (yxor_2__state == 2'b01);
  assign yxor_3___n__q0 = n;
  assign yxor_3__ap_start_global__q0 = ap_start__q0;
  assign yxor_3__is_done__q0 = (yxor_3__state == 2'b10);
  assign yxor_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_3__state <= 2'b00;
    end else begin
      if(yxor_3__state == 2'b00) begin
        if(yxor_3__ap_start_global__q0) begin
          yxor_3__state <= 2'b01;
        end
      end
      if(yxor_3__state == 2'b01) begin
        if(yxor_3__ap_ready) begin
          if(yxor_3__ap_done) begin
            yxor_3__state <= 2'b10;
          end else begin
            yxor_3__state <= 2'b11;
          end
        end
      end
      if(yxor_3__state == 2'b11) begin
        if(yxor_3__ap_done) begin
          yxor_3__state <= 2'b10;
        end
      end
      if(yxor_3__state == 2'b10) begin
        if(yxor_3__ap_done_global__q0) begin
          yxor_3__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_3__ap_start = (yxor_3__state == 2'b01);
  assign yxor_4___n__q0 = n;
  assign yxor_4__ap_start_global__q0 = ap_start__q0;
  assign yxor_4__is_done__q0 = (yxor_4__state == 2'b10);
  assign yxor_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_4__state <= 2'b00;
    end else begin
      if(yxor_4__state == 2'b00) begin
        if(yxor_4__ap_start_global__q0) begin
          yxor_4__state <= 2'b01;
        end
      end
      if(yxor_4__state == 2'b01) begin
        if(yxor_4__ap_ready) begin
          if(yxor_4__ap_done) begin
            yxor_4__state <= 2'b10;
          end else begin
            yxor_4__state <= 2'b11;
          end
        end
      end
      if(yxor_4__state == 2'b11) begin
        if(yxor_4__ap_done) begin
          yxor_4__state <= 2'b10;
        end
      end
      if(yxor_4__state == 2'b10) begin
        if(yxor_4__ap_done_global__q0) begin
          yxor_4__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_4__ap_start = (yxor_4__state == 2'b01);
  assign yxor_5___n__q0 = n;
  assign yxor_5__ap_start_global__q0 = ap_start__q0;
  assign yxor_5__is_done__q0 = (yxor_5__state == 2'b10);
  assign yxor_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_5__state <= 2'b00;
    end else begin
      if(yxor_5__state == 2'b00) begin
        if(yxor_5__ap_start_global__q0) begin
          yxor_5__state <= 2'b01;
        end
      end
      if(yxor_5__state == 2'b01) begin
        if(yxor_5__ap_ready) begin
          if(yxor_5__ap_done) begin
            yxor_5__state <= 2'b10;
          end else begin
            yxor_5__state <= 2'b11;
          end
        end
      end
      if(yxor_5__state == 2'b11) begin
        if(yxor_5__ap_done) begin
          yxor_5__state <= 2'b10;
        end
      end
      if(yxor_5__state == 2'b10) begin
        if(yxor_5__ap_done_global__q0) begin
          yxor_5__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_5__ap_start = (yxor_5__state == 2'b01);
  assign yxor_6___n__q0 = n;
  assign yxor_6__ap_start_global__q0 = ap_start__q0;
  assign yxor_6__is_done__q0 = (yxor_6__state == 2'b10);
  assign yxor_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_6__state <= 2'b00;
    end else begin
      if(yxor_6__state == 2'b00) begin
        if(yxor_6__ap_start_global__q0) begin
          yxor_6__state <= 2'b01;
        end
      end
      if(yxor_6__state == 2'b01) begin
        if(yxor_6__ap_ready) begin
          if(yxor_6__ap_done) begin
            yxor_6__state <= 2'b10;
          end else begin
            yxor_6__state <= 2'b11;
          end
        end
      end
      if(yxor_6__state == 2'b11) begin
        if(yxor_6__ap_done) begin
          yxor_6__state <= 2'b10;
        end
      end
      if(yxor_6__state == 2'b10) begin
        if(yxor_6__ap_done_global__q0) begin
          yxor_6__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_6__ap_start = (yxor_6__state == 2'b01);
  assign yxor_7___n__q0 = n;
  assign yxor_7__ap_start_global__q0 = ap_start__q0;
  assign yxor_7__is_done__q0 = (yxor_7__state == 2'b10);
  assign yxor_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_7__state <= 2'b00;
    end else begin
      if(yxor_7__state == 2'b00) begin
        if(yxor_7__ap_start_global__q0) begin
          yxor_7__state <= 2'b01;
        end
      end
      if(yxor_7__state == 2'b01) begin
        if(yxor_7__ap_ready) begin
          if(yxor_7__ap_done) begin
            yxor_7__state <= 2'b10;
          end else begin
            yxor_7__state <= 2'b11;
          end
        end
      end
      if(yxor_7__state == 2'b11) begin
        if(yxor_7__ap_done) begin
          yxor_7__state <= 2'b10;
        end
      end
      if(yxor_7__state == 2'b10) begin
        if(yxor_7__ap_done_global__q0) begin
          yxor_7__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_7__ap_start = (yxor_7__state == 2'b01);
  assign yxor_8___n__q0 = n;
  assign yxor_8__ap_start_global__q0 = ap_start__q0;
  assign yxor_8__is_done__q0 = (yxor_8__state == 2'b10);
  assign yxor_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_8__state <= 2'b00;
    end else begin
      if(yxor_8__state == 2'b00) begin
        if(yxor_8__ap_start_global__q0) begin
          yxor_8__state <= 2'b01;
        end
      end
      if(yxor_8__state == 2'b01) begin
        if(yxor_8__ap_ready) begin
          if(yxor_8__ap_done) begin
            yxor_8__state <= 2'b10;
          end else begin
            yxor_8__state <= 2'b11;
          end
        end
      end
      if(yxor_8__state == 2'b11) begin
        if(yxor_8__ap_done) begin
          yxor_8__state <= 2'b10;
        end
      end
      if(yxor_8__state == 2'b10) begin
        if(yxor_8__ap_done_global__q0) begin
          yxor_8__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_8__ap_start = (yxor_8__state == 2'b01);
  assign yxor_9___n__q0 = n;
  assign yxor_9__ap_start_global__q0 = ap_start__q0;
  assign yxor_9__is_done__q0 = (yxor_9__state == 2'b10);
  assign yxor_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_9__state <= 2'b00;
    end else begin
      if(yxor_9__state == 2'b00) begin
        if(yxor_9__ap_start_global__q0) begin
          yxor_9__state <= 2'b01;
        end
      end
      if(yxor_9__state == 2'b01) begin
        if(yxor_9__ap_ready) begin
          if(yxor_9__ap_done) begin
            yxor_9__state <= 2'b10;
          end else begin
            yxor_9__state <= 2'b11;
          end
        end
      end
      if(yxor_9__state == 2'b11) begin
        if(yxor_9__ap_done) begin
          yxor_9__state <= 2'b10;
        end
      end
      if(yxor_9__state == 2'b10) begin
        if(yxor_9__ap_done_global__q0) begin
          yxor_9__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_9__ap_start = (yxor_9__state == 2'b01);
  assign yxor_10___n__q0 = n;
  assign yxor_10__ap_start_global__q0 = ap_start__q0;
  assign yxor_10__is_done__q0 = (yxor_10__state == 2'b10);
  assign yxor_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_10__state <= 2'b00;
    end else begin
      if(yxor_10__state == 2'b00) begin
        if(yxor_10__ap_start_global__q0) begin
          yxor_10__state <= 2'b01;
        end
      end
      if(yxor_10__state == 2'b01) begin
        if(yxor_10__ap_ready) begin
          if(yxor_10__ap_done) begin
            yxor_10__state <= 2'b10;
          end else begin
            yxor_10__state <= 2'b11;
          end
        end
      end
      if(yxor_10__state == 2'b11) begin
        if(yxor_10__ap_done) begin
          yxor_10__state <= 2'b10;
        end
      end
      if(yxor_10__state == 2'b10) begin
        if(yxor_10__ap_done_global__q0) begin
          yxor_10__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_10__ap_start = (yxor_10__state == 2'b01);
  assign yxor_11___n__q0 = n;
  assign yxor_11__ap_start_global__q0 = ap_start__q0;
  assign yxor_11__is_done__q0 = (yxor_11__state == 2'b10);
  assign yxor_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_11__state <= 2'b00;
    end else begin
      if(yxor_11__state == 2'b00) begin
        if(yxor_11__ap_start_global__q0) begin
          yxor_11__state <= 2'b01;
        end
      end
      if(yxor_11__state == 2'b01) begin
        if(yxor_11__ap_ready) begin
          if(yxor_11__ap_done) begin
            yxor_11__state <= 2'b10;
          end else begin
            yxor_11__state <= 2'b11;
          end
        end
      end
      if(yxor_11__state == 2'b11) begin
        if(yxor_11__ap_done) begin
          yxor_11__state <= 2'b10;
        end
      end
      if(yxor_11__state == 2'b10) begin
        if(yxor_11__ap_done_global__q0) begin
          yxor_11__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_11__ap_start = (yxor_11__state == 2'b01);
  assign yxor_12___n__q0 = n;
  assign yxor_12__ap_start_global__q0 = ap_start__q0;
  assign yxor_12__is_done__q0 = (yxor_12__state == 2'b10);
  assign yxor_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_12__state <= 2'b00;
    end else begin
      if(yxor_12__state == 2'b00) begin
        if(yxor_12__ap_start_global__q0) begin
          yxor_12__state <= 2'b01;
        end
      end
      if(yxor_12__state == 2'b01) begin
        if(yxor_12__ap_ready) begin
          if(yxor_12__ap_done) begin
            yxor_12__state <= 2'b10;
          end else begin
            yxor_12__state <= 2'b11;
          end
        end
      end
      if(yxor_12__state == 2'b11) begin
        if(yxor_12__ap_done) begin
          yxor_12__state <= 2'b10;
        end
      end
      if(yxor_12__state == 2'b10) begin
        if(yxor_12__ap_done_global__q0) begin
          yxor_12__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_12__ap_start = (yxor_12__state == 2'b01);
  assign yxor_13___n__q0 = n;
  assign yxor_13__ap_start_global__q0 = ap_start__q0;
  assign yxor_13__is_done__q0 = (yxor_13__state == 2'b10);
  assign yxor_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_13__state <= 2'b00;
    end else begin
      if(yxor_13__state == 2'b00) begin
        if(yxor_13__ap_start_global__q0) begin
          yxor_13__state <= 2'b01;
        end
      end
      if(yxor_13__state == 2'b01) begin
        if(yxor_13__ap_ready) begin
          if(yxor_13__ap_done) begin
            yxor_13__state <= 2'b10;
          end else begin
            yxor_13__state <= 2'b11;
          end
        end
      end
      if(yxor_13__state == 2'b11) begin
        if(yxor_13__ap_done) begin
          yxor_13__state <= 2'b10;
        end
      end
      if(yxor_13__state == 2'b10) begin
        if(yxor_13__ap_done_global__q0) begin
          yxor_13__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_13__ap_start = (yxor_13__state == 2'b01);
  assign yxor_14___n__q0 = n;
  assign yxor_14__ap_start_global__q0 = ap_start__q0;
  assign yxor_14__is_done__q0 = (yxor_14__state == 2'b10);
  assign yxor_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_14__state <= 2'b00;
    end else begin
      if(yxor_14__state == 2'b00) begin
        if(yxor_14__ap_start_global__q0) begin
          yxor_14__state <= 2'b01;
        end
      end
      if(yxor_14__state == 2'b01) begin
        if(yxor_14__ap_ready) begin
          if(yxor_14__ap_done) begin
            yxor_14__state <= 2'b10;
          end else begin
            yxor_14__state <= 2'b11;
          end
        end
      end
      if(yxor_14__state == 2'b11) begin
        if(yxor_14__ap_done) begin
          yxor_14__state <= 2'b10;
        end
      end
      if(yxor_14__state == 2'b10) begin
        if(yxor_14__ap_done_global__q0) begin
          yxor_14__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_14__ap_start = (yxor_14__state == 2'b01);
  assign yxor_15___n__q0 = n;
  assign yxor_15__ap_start_global__q0 = ap_start__q0;
  assign yxor_15__is_done__q0 = (yxor_15__state == 2'b10);
  assign yxor_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_15__state <= 2'b00;
    end else begin
      if(yxor_15__state == 2'b00) begin
        if(yxor_15__ap_start_global__q0) begin
          yxor_15__state <= 2'b01;
        end
      end
      if(yxor_15__state == 2'b01) begin
        if(yxor_15__ap_ready) begin
          if(yxor_15__ap_done) begin
            yxor_15__state <= 2'b10;
          end else begin
            yxor_15__state <= 2'b11;
          end
        end
      end
      if(yxor_15__state == 2'b11) begin
        if(yxor_15__ap_done) begin
          yxor_15__state <= 2'b10;
        end
      end
      if(yxor_15__state == 2'b10) begin
        if(yxor_15__ap_done_global__q0) begin
          yxor_15__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_15__ap_start = (yxor_15__state == 2'b01);
  assign yxor_16___n__q0 = n;
  assign yxor_16__ap_start_global__q0 = ap_start__q0;
  assign yxor_16__is_done__q0 = (yxor_16__state == 2'b10);
  assign yxor_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_16__state <= 2'b00;
    end else begin
      if(yxor_16__state == 2'b00) begin
        if(yxor_16__ap_start_global__q0) begin
          yxor_16__state <= 2'b01;
        end
      end
      if(yxor_16__state == 2'b01) begin
        if(yxor_16__ap_ready) begin
          if(yxor_16__ap_done) begin
            yxor_16__state <= 2'b10;
          end else begin
            yxor_16__state <= 2'b11;
          end
        end
      end
      if(yxor_16__state == 2'b11) begin
        if(yxor_16__ap_done) begin
          yxor_16__state <= 2'b10;
        end
      end
      if(yxor_16__state == 2'b10) begin
        if(yxor_16__ap_done_global__q0) begin
          yxor_16__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_16__ap_start = (yxor_16__state == 2'b01);
  assign yxor_17___n__q0 = n;
  assign yxor_17__ap_start_global__q0 = ap_start__q0;
  assign yxor_17__is_done__q0 = (yxor_17__state == 2'b10);
  assign yxor_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_17__state <= 2'b00;
    end else begin
      if(yxor_17__state == 2'b00) begin
        if(yxor_17__ap_start_global__q0) begin
          yxor_17__state <= 2'b01;
        end
      end
      if(yxor_17__state == 2'b01) begin
        if(yxor_17__ap_ready) begin
          if(yxor_17__ap_done) begin
            yxor_17__state <= 2'b10;
          end else begin
            yxor_17__state <= 2'b11;
          end
        end
      end
      if(yxor_17__state == 2'b11) begin
        if(yxor_17__ap_done) begin
          yxor_17__state <= 2'b10;
        end
      end
      if(yxor_17__state == 2'b10) begin
        if(yxor_17__ap_done_global__q0) begin
          yxor_17__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_17__ap_start = (yxor_17__state == 2'b01);
  assign yxor_18___n__q0 = n;
  assign yxor_18__ap_start_global__q0 = ap_start__q0;
  assign yxor_18__is_done__q0 = (yxor_18__state == 2'b10);
  assign yxor_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_18__state <= 2'b00;
    end else begin
      if(yxor_18__state == 2'b00) begin
        if(yxor_18__ap_start_global__q0) begin
          yxor_18__state <= 2'b01;
        end
      end
      if(yxor_18__state == 2'b01) begin
        if(yxor_18__ap_ready) begin
          if(yxor_18__ap_done) begin
            yxor_18__state <= 2'b10;
          end else begin
            yxor_18__state <= 2'b11;
          end
        end
      end
      if(yxor_18__state == 2'b11) begin
        if(yxor_18__ap_done) begin
          yxor_18__state <= 2'b10;
        end
      end
      if(yxor_18__state == 2'b10) begin
        if(yxor_18__ap_done_global__q0) begin
          yxor_18__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_18__ap_start = (yxor_18__state == 2'b01);
  assign yxor_19___n__q0 = n;
  assign yxor_19__ap_start_global__q0 = ap_start__q0;
  assign yxor_19__is_done__q0 = (yxor_19__state == 2'b10);
  assign yxor_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_19__state <= 2'b00;
    end else begin
      if(yxor_19__state == 2'b00) begin
        if(yxor_19__ap_start_global__q0) begin
          yxor_19__state <= 2'b01;
        end
      end
      if(yxor_19__state == 2'b01) begin
        if(yxor_19__ap_ready) begin
          if(yxor_19__ap_done) begin
            yxor_19__state <= 2'b10;
          end else begin
            yxor_19__state <= 2'b11;
          end
        end
      end
      if(yxor_19__state == 2'b11) begin
        if(yxor_19__ap_done) begin
          yxor_19__state <= 2'b10;
        end
      end
      if(yxor_19__state == 2'b10) begin
        if(yxor_19__ap_done_global__q0) begin
          yxor_19__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_19__ap_start = (yxor_19__state == 2'b01);
  assign yxor_20___n__q0 = n;
  assign yxor_20__ap_start_global__q0 = ap_start__q0;
  assign yxor_20__is_done__q0 = (yxor_20__state == 2'b10);
  assign yxor_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_20__state <= 2'b00;
    end else begin
      if(yxor_20__state == 2'b00) begin
        if(yxor_20__ap_start_global__q0) begin
          yxor_20__state <= 2'b01;
        end
      end
      if(yxor_20__state == 2'b01) begin
        if(yxor_20__ap_ready) begin
          if(yxor_20__ap_done) begin
            yxor_20__state <= 2'b10;
          end else begin
            yxor_20__state <= 2'b11;
          end
        end
      end
      if(yxor_20__state == 2'b11) begin
        if(yxor_20__ap_done) begin
          yxor_20__state <= 2'b10;
        end
      end
      if(yxor_20__state == 2'b10) begin
        if(yxor_20__ap_done_global__q0) begin
          yxor_20__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_20__ap_start = (yxor_20__state == 2'b01);
  assign yxor_21___n__q0 = n;
  assign yxor_21__ap_start_global__q0 = ap_start__q0;
  assign yxor_21__is_done__q0 = (yxor_21__state == 2'b10);
  assign yxor_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_21__state <= 2'b00;
    end else begin
      if(yxor_21__state == 2'b00) begin
        if(yxor_21__ap_start_global__q0) begin
          yxor_21__state <= 2'b01;
        end
      end
      if(yxor_21__state == 2'b01) begin
        if(yxor_21__ap_ready) begin
          if(yxor_21__ap_done) begin
            yxor_21__state <= 2'b10;
          end else begin
            yxor_21__state <= 2'b11;
          end
        end
      end
      if(yxor_21__state == 2'b11) begin
        if(yxor_21__ap_done) begin
          yxor_21__state <= 2'b10;
        end
      end
      if(yxor_21__state == 2'b10) begin
        if(yxor_21__ap_done_global__q0) begin
          yxor_21__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_21__ap_start = (yxor_21__state == 2'b01);
  assign yxor_22___n__q0 = n;
  assign yxor_22__ap_start_global__q0 = ap_start__q0;
  assign yxor_22__is_done__q0 = (yxor_22__state == 2'b10);
  assign yxor_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_22__state <= 2'b00;
    end else begin
      if(yxor_22__state == 2'b00) begin
        if(yxor_22__ap_start_global__q0) begin
          yxor_22__state <= 2'b01;
        end
      end
      if(yxor_22__state == 2'b01) begin
        if(yxor_22__ap_ready) begin
          if(yxor_22__ap_done) begin
            yxor_22__state <= 2'b10;
          end else begin
            yxor_22__state <= 2'b11;
          end
        end
      end
      if(yxor_22__state == 2'b11) begin
        if(yxor_22__ap_done) begin
          yxor_22__state <= 2'b10;
        end
      end
      if(yxor_22__state == 2'b10) begin
        if(yxor_22__ap_done_global__q0) begin
          yxor_22__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_22__ap_start = (yxor_22__state == 2'b01);
  assign yxor_23___n__q0 = n;
  assign yxor_23__ap_start_global__q0 = ap_start__q0;
  assign yxor_23__is_done__q0 = (yxor_23__state == 2'b10);
  assign yxor_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_23__state <= 2'b00;
    end else begin
      if(yxor_23__state == 2'b00) begin
        if(yxor_23__ap_start_global__q0) begin
          yxor_23__state <= 2'b01;
        end
      end
      if(yxor_23__state == 2'b01) begin
        if(yxor_23__ap_ready) begin
          if(yxor_23__ap_done) begin
            yxor_23__state <= 2'b10;
          end else begin
            yxor_23__state <= 2'b11;
          end
        end
      end
      if(yxor_23__state == 2'b11) begin
        if(yxor_23__ap_done) begin
          yxor_23__state <= 2'b10;
        end
      end
      if(yxor_23__state == 2'b10) begin
        if(yxor_23__ap_done_global__q0) begin
          yxor_23__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_23__ap_start = (yxor_23__state == 2'b01);
  assign yxor_24___n__q0 = n;
  assign yxor_24__ap_start_global__q0 = ap_start__q0;
  assign yxor_24__is_done__q0 = (yxor_24__state == 2'b10);
  assign yxor_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_24__state <= 2'b00;
    end else begin
      if(yxor_24__state == 2'b00) begin
        if(yxor_24__ap_start_global__q0) begin
          yxor_24__state <= 2'b01;
        end
      end
      if(yxor_24__state == 2'b01) begin
        if(yxor_24__ap_ready) begin
          if(yxor_24__ap_done) begin
            yxor_24__state <= 2'b10;
          end else begin
            yxor_24__state <= 2'b11;
          end
        end
      end
      if(yxor_24__state == 2'b11) begin
        if(yxor_24__ap_done) begin
          yxor_24__state <= 2'b10;
        end
      end
      if(yxor_24__state == 2'b10) begin
        if(yxor_24__ap_done_global__q0) begin
          yxor_24__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_24__ap_start = (yxor_24__state == 2'b01);
  assign yxor_25___n__q0 = n;
  assign yxor_25__ap_start_global__q0 = ap_start__q0;
  assign yxor_25__is_done__q0 = (yxor_25__state == 2'b10);
  assign yxor_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_25__state <= 2'b00;
    end else begin
      if(yxor_25__state == 2'b00) begin
        if(yxor_25__ap_start_global__q0) begin
          yxor_25__state <= 2'b01;
        end
      end
      if(yxor_25__state == 2'b01) begin
        if(yxor_25__ap_ready) begin
          if(yxor_25__ap_done) begin
            yxor_25__state <= 2'b10;
          end else begin
            yxor_25__state <= 2'b11;
          end
        end
      end
      if(yxor_25__state == 2'b11) begin
        if(yxor_25__ap_done) begin
          yxor_25__state <= 2'b10;
        end
      end
      if(yxor_25__state == 2'b10) begin
        if(yxor_25__ap_done_global__q0) begin
          yxor_25__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_25__ap_start = (yxor_25__state == 2'b01);
  assign yxor_26___n__q0 = n;
  assign yxor_26__ap_start_global__q0 = ap_start__q0;
  assign yxor_26__is_done__q0 = (yxor_26__state == 2'b10);
  assign yxor_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_26__state <= 2'b00;
    end else begin
      if(yxor_26__state == 2'b00) begin
        if(yxor_26__ap_start_global__q0) begin
          yxor_26__state <= 2'b01;
        end
      end
      if(yxor_26__state == 2'b01) begin
        if(yxor_26__ap_ready) begin
          if(yxor_26__ap_done) begin
            yxor_26__state <= 2'b10;
          end else begin
            yxor_26__state <= 2'b11;
          end
        end
      end
      if(yxor_26__state == 2'b11) begin
        if(yxor_26__ap_done) begin
          yxor_26__state <= 2'b10;
        end
      end
      if(yxor_26__state == 2'b10) begin
        if(yxor_26__ap_done_global__q0) begin
          yxor_26__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_26__ap_start = (yxor_26__state == 2'b01);
  assign yxor_27___n__q0 = n;
  assign yxor_27__ap_start_global__q0 = ap_start__q0;
  assign yxor_27__is_done__q0 = (yxor_27__state == 2'b10);
  assign yxor_27__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_27__state <= 2'b00;
    end else begin
      if(yxor_27__state == 2'b00) begin
        if(yxor_27__ap_start_global__q0) begin
          yxor_27__state <= 2'b01;
        end
      end
      if(yxor_27__state == 2'b01) begin
        if(yxor_27__ap_ready) begin
          if(yxor_27__ap_done) begin
            yxor_27__state <= 2'b10;
          end else begin
            yxor_27__state <= 2'b11;
          end
        end
      end
      if(yxor_27__state == 2'b11) begin
        if(yxor_27__ap_done) begin
          yxor_27__state <= 2'b10;
        end
      end
      if(yxor_27__state == 2'b10) begin
        if(yxor_27__ap_done_global__q0) begin
          yxor_27__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_27__ap_start = (yxor_27__state == 2'b01);
  assign yxor_28___n__q0 = n;
  assign yxor_28__ap_start_global__q0 = ap_start__q0;
  assign yxor_28__is_done__q0 = (yxor_28__state == 2'b10);
  assign yxor_28__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yxor_28__state <= 2'b00;
    end else begin
      if(yxor_28__state == 2'b00) begin
        if(yxor_28__ap_start_global__q0) begin
          yxor_28__state <= 2'b01;
        end
      end
      if(yxor_28__state == 2'b01) begin
        if(yxor_28__ap_ready) begin
          if(yxor_28__ap_done) begin
            yxor_28__state <= 2'b10;
          end else begin
            yxor_28__state <= 2'b11;
          end
        end
      end
      if(yxor_28__state == 2'b11) begin
        if(yxor_28__ap_done) begin
          yxor_28__state <= 2'b10;
        end
      end
      if(yxor_28__state == 2'b10) begin
        if(yxor_28__ap_done_global__q0) begin
          yxor_28__state <= 2'b00;
        end
      end
    end
  end

  assign yxor_28__ap_start = (yxor_28__state == 2'b01);

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      tapa_state <= 2'b00;
    end else begin
      case(tapa_state)
        2'b00: begin
          if(ap_start__q0) begin
            tapa_state <= 2'b01;
          end
        end
        2'b01: begin
          if(Mmap2Stream_0__is_done__q0 && Mmap2Stream_1__is_done__q0 && Mmap2Stream_2__is_done__q0 && Mmap2Stream_3__is_done__q0 && Mmap2Stream_4__is_done__q0 && Mmap2Stream_5__is_done__q0 && Mmap2Stream_6__is_done__q0 && Mmap2Stream_7__is_done__q0 && Mmap2Stream_8__is_done__q0 && Mmap2Stream_9__is_done__q0 && Mmap2Stream_10__is_done__q0 && Mmap2Stream_11__is_done__q0 && Mmap2Stream_12__is_done__q0 && Mmap2Stream_13__is_done__q0 && Mmap2Stream_14__is_done__q0 && Mmap2Stream_15__is_done__q0 && Mmap2Stream_16__is_done__q0 && Mmap2Stream_17__is_done__q0 && Mmap2Stream_18__is_done__q0 && Mmap2Stream_19__is_done__q0 && Mmap2Stream_20__is_done__q0 && Mmap2Stream_21__is_done__q0 && Mmap2Stream_22__is_done__q0 && Mmap2Stream_23__is_done__q0 && Mmap2Stream_24__is_done__q0 && Mmap2Stream_25__is_done__q0 && Mmap2Stream_26__is_done__q0 && Mmap2Stream_27__is_done__q0 && Mmap2Stream_28__is_done__q0 && Mmap2Stream_29__is_done__q0 && Stream2Mmap_0__is_done__q0 && yxor_0__is_done__q0 && yxor_1__is_done__q0 && yxor_2__is_done__q0 && yxor_3__is_done__q0 && yxor_4__is_done__q0 && yxor_5__is_done__q0 && yxor_6__is_done__q0 && yxor_7__is_done__q0 && yxor_8__is_done__q0 && yxor_9__is_done__q0 && yxor_10__is_done__q0 && yxor_11__is_done__q0 && yxor_12__is_done__q0 && yxor_13__is_done__q0 && yxor_14__is_done__q0 && yxor_15__is_done__q0 && yxor_16__is_done__q0 && yxor_17__is_done__q0 && yxor_18__is_done__q0 && yxor_19__is_done__q0 && yxor_20__is_done__q0 && yxor_21__is_done__q0 && yxor_22__is_done__q0 && yxor_23__is_done__q0 && yxor_24__is_done__q0 && yxor_25__is_done__q0 && yxor_26__is_done__q0 && yxor_27__is_done__q0 && yxor_28__is_done__q0) begin
            tapa_state <= 2'b10;
          end
        end
        2'b10: begin
          tapa_state <= 2'b00;
          countdown <= 1'd0;
        end
        2'b11: begin
          if(countdown == 1'd0) begin
            tapa_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end
      endcase
    end
  end

  assign ap_idle = (tapa_state == 2'b00);
  assign ap_done = ap_done__q0;
  assign ap_ready = ap_done__q0;
  assign ap_start__q0 = ap_start;
  assign ap_done__q0 = (tapa_state == 2'b10);

endmodule
