(* DONT_TOUCH = "yes" *)
module gnd_driver(
    output dout
    );

    assign dout = 1'b0;

endmodule
